ELF              �4   �#     4    (           � �� �          � DD�   8'           � DD             U���D  �?h ]�             S���H�Y��ɉXQQRP�� ����[�f�f�f�f�f�f�f��=�E u��E�=�E u��E�=�E u��E�=�E u��E�=xE u�xE�=pE u�pE�=hE u�hE�=`E u�`E�=XE u�XE�=PE u�PE�=HE u�HE�=@E u�@E��f�f�f�f�f�f�f���h`Dh�Dh�'裲 ��h`Dh�Dh�'茲 ���蒲 ���f�f�f���D-�D��v�    ��tU���h�D�Ѓ���Ð�t& ��D-�D���������t�    ��tU���Ph�D�҃���Ít& ��'    �= E uhU��S�4D��0D���E����9�s��    ���E��0D�E9�r��C���� -��t��h��	�]� ��� E�]���Í�    ��'    U�`*�����t��hEh��	�_� ���8D���u������t& ��'    �    ��t��P�҃���U��    ]ÍL$����q�U��SQ���   ��h���y� ����������   ��jj�  ����P�����P�A� ����h���������P��*  ����h��P��*  ���Ẽ������RP�p� �����E�P��  �����E�P�R	 ���   �������P�{ ���H  �   ��P�y� ���8E�8E��u^���E�P��j �����E�Ph���E�P��$ �����E�P�c  �����E�P�� �����E�P�j ���   ��   �8E�@�8E�@	 �8E� �8E�@ �  ��  �E�   �E��P�&  ���E��<� �E���u��u�貪 ���E�}�ua�E��E�E����E��E� ��P�ݩ ���Eܺ   �8E���u�RP�k� ���E؋E؉EȋE�P�E� Rj�U�RP覫 ��냉��a�Ã��E�P�� ����Ã������P�z ���؃�P赐 �Ã��E�P� ����Ã��E�P�i ���؃�P膐 �e�Y[]�a��U��S�����j`�M
  ����jd�@
  ������������u׃�j �m  ����h�   jd�0
  ����j �N  ����j jd�
  ����j�2  ����j`��	  �����E���j �  ����j`jd��	  ����j ��  ���E���Pj`�	  ����h�   �U  ����j��  ����j`�q	  ���E��}��tY���E�P�Eh �����E�Ph��E�P�]" �����E�P��  �����E�P�? �����E�P� h ����   ��h�   ��  ����j�;  ����j`��  ���E��}����   ���E�P�g �����E�PhD��E�P��! �����E�P�@  �����E�P� �����E�P�g ����^�Ã��E�P� ����Ã��E�P�ig ���؃�P�k� �Ã��E�P�] ����Ã��E�P�:g ���؃�P�<� �]���U���(�E�E�� E����t9��tI����   �E�!E�E����u� E ��   � E��   �E�"E� E�   �E�#E�!E�E��"E�E��#E�E��E���@��u�}� xy�E��U���f�� )�f�E��E��U���f�� )�f�E�8E����P�ҥ ���8E�U�f�P�8E�U�f�P�8Ef�U�f�P�8E�  �8E�@� E ���U����E�E��8E��	��P�o� ���8E�U�P
�8E�@ �8E�@	��U����E��� �} u4���jd�  ������������t�L�E�P��U������u��8�}u2���jd�^  ������������t��E�P��U������u���U����E�E��j �i�������h�   jd�,  ����j �J������E��Pj`�  ����U����}u3�}��  u*��h<E�dk ����h`Dh<Eh����� ����U�����h��  j��������U��U�E	�]�U��    ]�U��S�����E�P�Qd �����E�Ph���E�P�i �����E�P��  �����E�P�K �����E�P�,d ����ha�j�?� ����ha�j�-� ���/�Ã��E�P� ����Ã��E�P��c ���؃�P�� �]���U���(�E�E��c��j`�  ���E��E��� �����E��}� t�E���P��������E���P�V������0E�4E���� �0E�4E��jd�H  ���E��E����������y�����U����}u3�}��  u*��h=E�i ����h`Dh=Eh���6� ����U�����h��  j��������U��    ]�U����}u3�}��  u*��h>E�Ai ����h`Dh>Eh���ѧ ����U�����h��  j��������U��    ]�U��S��  ��h   �  ���E���u��F� ����h��Z� �����u��� ����P�v  ����jh#��� ���P�#� ���ܡ �Ã�h+��� �����P�2!  ����SP��&  ����h.�P�!  �����uP�6  ����h �P�d  �����u�躣 �����u��8  ������ ���P��� ������ ���P�� ����Ã��� ���P�n� ���؃�P�P� �]���U����}u3�}��  u*��h?E�g ����h`Dh?Eh���9� ����U�����h��  j��������U��    ]�U��S���E�E�]���u�{� ����SP�(   ���]���U����E�E�E��P�u�   ����U������u�y0 ���E�E���E��E���P�  ���E��u�u�u��u��( �����u��|� �����u���  ���ÐU��    ]�U��S���E�    ��E��E��P�u�% ��� ����P�U� ��������uσ��u��� ���E���m��E�����P�u��  ��� ����P�� ��������űE�;E�7���E�P�\_ �����E�PhA��u�u �����E�P�V_ ���:�E�+E���U�EQR�uP�� ����Ã��E�P�%_ ���؃�P�'� �E�]��� �U����Ef�E��E���E��E��ÐU����U�Ef�U��E��U��E����U����Ef�E��E��f�f�E��E��ÐU����U�Ef�U�f�E��U��E�f���U����Ef�E��E���E��E���U����Ef�E��U��E���f�f�f�f�f�f���t� f�f�f�f�f��WV��S1�1ɍ�&    ���P��Ӄ����	ބ�x��w��@t	�������	։7[^_�WV��S�ωӃ���D$�R�P����t
�D$� �D$j��T$RSV�P����t�T$���[^_�f�f��UW��VS�΃�,<P�T$��   ����<��   ���$���f���Y��t����p<Et$����y��D$@���,��[^_]Ð��Y�Ή���'    ��Y뽐��&    �T$��������T$��뢍�    ��'    1҉�1ɉՐ��&    ���S��Ѓ�����	ń�x���g���f���Y�Z�����t& �% �t& ��'    ���D$@�����^���,��[^_]�f�f��S���X���ts�ك���tYv7��t6���ڀ�u8�H��ыP�Í\$S�����D$��([Í�&    ��u�����͐�t& �'% �t& ��'    ���벍v ��'    1��f�f�f�f�f�f�UW��VS�ǃ��t$0�L$��p���&    1�1ɍ�    ��    ���F��Ã����	ڄ�x��t�������L$��������t���[^_]Ã�1�[^_]�f�f�f�f�f�f����<�t)��p< tRv0<@t<<Pt<0u,��R�K ����Ít& 1���Ív ��'    ��t�<t��/$ �v ��R�~ ����Ã�R� �����UW��VS1��Ճ����L$t��W�~ ���\$�u��U �����   ������M����S����R������������V�t$<��F��   1�1ɍ�    ��'    ���Z��؃�����	Ǆ�x�D$׉x�B��t$1�1ɈV�����������������X��ڃ����	ׄ�x�t$ǉ~��[^_]Ð��&    �|$�G�^����t& �D$�@    �f��UW�   VS��\�|$p�L$x�\$|�D$$    �D$(    t��\[^_]Í�    ��'    �� �Լ�D$�Ӽ����� ��   �|$t��8D$��   ��$�   �X�@��D$��$�   �p����  �D$t�  ����  ����$�   j ��$�   �| ��Sj��$�   �| XZV��$�   �| ���   ��\[^_]Ð�t& ���D$�|$t��8D$�b�������$�   �g| �D$������  �T$��$�   �L$8�������D$L��$�   �1������D$H�D$0P��$�   ��{ ���ƃ|$(�� ;\$H��   �|$,�l$M1҉���������ى�W��������\$]�Ń�1҉����������D$<P�������\$]�Ń�1҉���������D$@1�P���s�������1ɍ�    ��    ���S��Ѓ�����	ń�x�D$8D$,9���   1��   1�1��D$t��   ����   �|$ �   �������$�   �L$�W�T$$�_�O��w�W�������&    �D$tuy����$�   �  �v ��'    ��t[��������. ��&    ��'    �D$tuـ|$ u҃������뮍�&    D$09�r';\$H������0�������'    �+. �   �����D$4��t�D$<����0  �D$H���D(���t҅��"  �D$t�D$@	���D$u3�|$ �D$�	u$��$�   ��$�   �� �t�GЉD$$�@��D$�D$ �׉t$f��T$0���5����T$4���*����T$0�� tej�L$�\$��������!�:D$��   ��T$D1�1ɍ�&    ���Z��؃�����	ń�x������uA�D$4����   �<�|����D$��D$8�L�����t�l$��tЋT$�L$$�������t����t$�\$0�   �������������   ������T$��$�   �L$8�u����D$L��$�   ������D$@�D$L��$�   �������$�   �G��������R�L$4�T$ �D$H�;��������,����|$ ���t$�$���1۸   �E�����P��& �5, f�f��U��WVS��H�]S��& �C��s�{܉EċC�E�X�s��, ��P�& �u& � ���@0�XPt��UčM�1��������S��E�V����������t�K  ����& ��& ��S�{ ���E�1�V��	�c�������t#��j�b, ��� �	h0�h�	P�   ��W� + U����u�- ���Ã�t	��P�/{ ��P����f�f�f�S���|$�D$w6��h�u*�PԍX ��t	��S�҃��\$��[�Z, �v ��'    ��[Ã��p��* S���\$�c% �@�D$�C�   �� �CЋD$�C��+ �C���* � ++C�C܃��CCUNG�C �S�Zx �$�2% �}* f�f�f�f�f�f��S����$ ��@��t4�J0�Z4�� �Լ�Ӽ����� v"�     �Z0��S��z �$��$ ���$* ��w��Z��f�f�f�f�f�S���\$��t4��S�$ ��S �Լ�Ҽ������� w��w���s��) �v ��) f�f�f�f�f���D$�f�f�f�f�f��D$� L��@�	���D$�� �v �D$�A�D$�ѐS���\$�C�L��C�	P�� �\$ ��[�������t& �D$�A�D$����T$�D$�
�A�R��T$�D$�T$�� f�f�f�f�f��U��WVS���]�sV�� �Ct    �Cx �Cy �C|    ǃ�       ǃ�       ǃ�       �L��C`�XZ�uV�� ���e�[^_]Éǃ��C�	V�� �<$�zx f�f�f�f�f��L$�D$���R�I��f�f�f�f�f��D$��f�f�f�f�f�S���\$��P��R�T$$����[�f�f��S���\$��P��R�T$$����[�f�f��VS���\$�t$��@�Dx�V�t$P�R0��9�t(�X�C�\$���D$��[^鋜 �t& ��'    ��[^�f�f�f�f�f�U��S���]��@�Dx��t���P�R�����t�؋]��Ð����P�ڋB��PR�)� �؃��]��Ã�u ��P�" ���X�K�Ct-�������P��! ����H�كI�Au�H" 뎉��
���������3" ��S��v ���#" ��S��v f�f�f�f�f�U��VS���u�]�������C�����H���At�e���[^]� ��    ��'    �Ax�M���jjj j PQ�R�E����E��C�E�C�e���[^]� ��u ��P�
! ���p�N�Ft.�������P��  ���p�N�Fu�S! �f������
���������;! ��S��u ���+! ��S��u f�U��WVS��,�]��x���Gt�e��[^_]Í�    ��'    �Gx�U���M�u�8jVQRP�EЉU܉M��u�P�W�E�#Eԃ����u�����P�ڋB��PR�4� ��똃�u ��P�  ���X�K�Ct0�������P�� ����H�كI�Au�X  �L������
���������@  ��S��t ���0  ��S��t f�f�f��U��WVS���]�u�}��H���At�e��[^_]Í�&    �Ax�M܃��j�uWVPQ�R�E�#E������uʋ���P�ڋB��PR�D� ��뮃�u ��P�! ���X�K�Ct0�������P� ����x�߃O�Gu�h �b������
���������P ��S�t ���@ ��S��s f�f�f���T$�D$�
�A�R��D$    �D$髝 f�f�f�f�f��U��WVS���]�sV��| �Ct    �Cx �Cy �C|    ǃ�       ǃ�       ǃ�       �L��C`�XZj V�@� ���e�[^_]Éǃ��C�	V�� �<$�;s f�f�f�f�f��VS���\$�t$��^� �H�ىȋIp��t�P��u&��Q�]������X�S�؅�u���[^Ív ���D$�T$��[^雗 f�f�f�f�f��VS���t$�F�B��@ ��t!�b ��u�Cx��t���P�R�����t��[^ËF���B�P��RP�8� ����[^�f�f�f�f�f�f�f��U��WVS�}���$�u�]VW���������|   �}� tv�E߃�P��@��txS�V ����u�����J��APQ�Ö ���U��X���C t!� ��u�Cx��t���P�R�����t�e��[^_]Ð�t& ��u��   랐�t& �E���B�P��RP�X� ���e��[^_]É���� ��W�����$�_q ��u ��P� ���p�N�Ft0�������P�� ����H��I�Au�X �#�����������������> �f�f�f�f�f�f�U��WVS�]���$�u�}VS�������}� t��@�Dx�P;Ps}���
�@�U��X���C t!�` ��u�Cx��t���P�R�����t�e��[^_]Ív ��'    �E���B�P��RP�(� ���e��[^_]Ít& ��'    �������WP�R4������p�������P��B��PR�ޔ ���Q�������*��u?��P� ���p�N�Ft�{���� ��S�����4$��o �����\�����P�s ����H��I�Au
�� ������0������� �f�f�f��U��WVS�}���$�u�]VW�7������}� t7����@�Dx�S�uP�R0��9�t����P��B��PR��� ���U��X���C t!�� ��u�Cx��t���P�R�����t�e��[^_]Í�    ��    �E���B�P��RP蘓 ���e��[^_]Ã�u ��P�m ���p�N�Ft0�6�����P�M ����H��I�Au-� �H����������� ��W�����$�Pn ������������ ��f�f�f�f�f�f�f��D$� �f�f�f�f�VS���t$��@�\|��tX�{ t$�C'��PV�����D$ ��[^�H������&    ��S�H ����P�
   ����t�j
S�҃�����- f�f�f�f�f�f����j �t$�������f�f�f�f�f�f�f������f�f�f�f�f��WVS�\$��p�ހ~u t�D$�Ft��[^_Í�&    ��'    �~|��t>� t�D$�Fu�Ft��[^_Ð��W��G ����@=��tՃ�j W�Ѓ����v f�f�f��D$��J���ʋL$	J�f�f�f�f�f���D$��J�T$���!Q�f�f�f�f�f��S�T$�D$��t2��
�   t1Ƀ�������Z�ËS��	ʉS[É���'    �@   ��f�f�f�f���D$�L$��R�L�f�f�f�f�f�f�f��D$�L$��R�L�f�f�f�f�f�f�f�U��WVS�E���4�]SP��������}� tK��@�<�w;u�}Љu�~{�O�ʉMԁ�   �� ���E��MԄ��h  �r����   �B    �E�B��@ ��t%�a ��u�Fx��t���P�R�������  �e��[^_]Í�&    �EЃ��@x��u�uP�R0��9E�ڋtP���B��PR�� �����P��p�����    ��'    �Bx����u�uP�R0��9Et����P�ڋB��PR迏 ���}� t���@�<�O���������u�+u�u �1  �Ot���Mԅ�������}��"�v ��'    �MԈ
�@����T����@�Dx�P;Pr܋��WP�R4�����uԋ�������+u�u �  �t���������ɉM��#��    ��'    ���
�@����}   �@�Dx�P;Prދ���u�P�R4�����uҋ���P�ڋB��PR賎 ����P�������t& �E���B�P��RP舎 ���e��[^_]Ít& ��'    �P���������    �G|���E���   �EԀx tY�@=�E��E��Gu�Gt��@������v ��'    �EЋx|��tw� tP�=�MЉ��At��Au�@�������v ���u���C �Eԃ�� �@=��uO�E� 닍�    ��'    ��W��C ����@=��u�    ��/�J� �E� RRj W�Љǃ��x���RRj �u��ЈEԃ��.�����u ��P�R ���X�K�Ct0������P�2 ����p�ރN�Fu0� ������������� �E���P�z����$�2h ������������b �ڃ� �D$(�D$j�D$P�t$,�������,Ð�� �D$(�D$j�D$P�t$,�������,Ð�� �D$(�D$j�D$P�t$,������,ÐVS���\$�t$��t��S� ��PSV�{���������[^Ë���P��B��PR�I� ������[^�f�f�f�f�f�f�f�VS���\$�t$��t��S�: ��PSV����������[^Ë���P��B��PR�� ������[^�f�f�f�f�f�f�f�VS���\$�t$��t��S�� ��PSV����������[^Ë���P��B��PR艋 ������[^�f�f�f�f�f�f�f�U��WVS�E���4�uVP�Z������}� tk��X�󋻀   ���N  �{u ��   �Ct�E̋Kx1҅ɉȋ���u�u�SRP�E�WP�Q���}� t����P��B��PR�� ���E�B��@ ��t!�� ��u�Cx��t���P�R�����tU�e��[^_]Ít& ��'    �C|���E���   �EȀx tY�H=�ȉM̈Ct��Cu�X���B�����    ��'    �E���B�P��RP�H� ���e��[^_]Ít& ��'    ���u��5@ �Eȃ��E�    � �P�    ����t���j �u����ȃ��M��n����� �	�� ���*��uB��P�� ���p�N�Ft"�����$ �E���P�����$��d �����g�����P�~ ����x���O�Gu
�� �����;������� �f������f�f�f�f�f���T$�L$��@�D��J��t��@t�ɉT$�L$����f��ɉT$�L$��������f�f�f�f�f��U��WVS�E���4�uVP��������}� tk��X�󋻀   ���N  �{u ��   �Ct�E̋Kx1҅ɉȋ���u�u�SRP�E�WP�Q���}� t����P��B��PR�y� ���E�B��@ ��t!�Q ��u�Cx��t���P�R�����tU�e��[^_]Ít& ��'    �C|���E���   �EȀx tY�H=�ȉM̈Ct��Cu�X���B�����    ��'    �E���B�P��RP�؇ ���e��[^_]Ít& ��'    ���u���= �Eȃ��E�    � �P�    ����t���j �u����ȃ��M��n����)� �	�"� ���*��uB��P�P ���p�N�Ft"����� �E���P�����$�`b �����������P� ����x���O�Gu
�u ������������d �f������f�f�f�f�f���D$�D$�����f������f�f�f�f�f��U��WVS��D�E�]�EčE�SP�������}� tz��x�ߋ��   ���X  �u ��   �Gt���E��yx�Uċ�E�    ���}ȍ}��Ẽ�R�u�Q�u��u�VW�P���}� t����P�ڋB��PR�$� ���E�B��@ ��t!�� ��u�Fx��t���P�R�����tP�e��[^_]Í�    �G|���E���   �EȀx tY�H=�ȉM��Gt��Gu�H���:�����    ��'    �E���B�P��RP舅 ���e��[^_]Ít& ��'    ���u��u; �Eȃ��E�    � �P�    ����t���j �u����ȃ��M��n������ �	��� ���*��uB��P�  ���X�K�Ct"������d �E���P�X����$�` ����������P�
 ����H�كI�Au
�% �����{������ �f��D$�D$�����f�U��WVS��D�E�u�U�EȍE�V�U�P�n������}� tk��X�󋻀   ���R  �{u ��   �Ct�EċKx1҅ɉȋ���u��u��u�SRP�E�WP�Q���}� t����P��B��PR��� ���E�B��@ ��t!��
 ��u�Cx��t���P�R�����tY�e��[^_]����������������C|���E���   �E��x tY�H=�ȉMĈCt��Cu�X���>�����    ��'    �E���B�P��RP�X� ���e��[^_]Ít& ��'    ���u��E9 �E����E�    � �P�    ����t���j �u����ȃ��M��n����� �	�� ���*��uB��P�� ���p�N�Ft"�����4	 �E���P�(����$��] �����w�����P� ����x���O�Gu
�� �����K������� �f������f�f�f�f�f��U��WVS��D�E�u�U�EȍE�V�U�P�>������}� tk��X�󋻀   ���R  �{u ��   �Ct�EċKx1҅ɉȋ���u��u��u�SRP�E�WP�Q���}� t����P��B��PR�́ ���E�B��@ ��t!� ��u�Cx��t���P�R�����tY�e��[^_]����������������C|���E���   �E��x tY�H=�ȉMĈCt��Cu�X���>�����    ��'    �E���B�P��RP�(� ���e��[^_]Ít& ��'    ���u��7 �E����E�    � �P�    ����t���j �u����ȃ��M��n����y� �	�r� ���*��uB��P� ���p�N�Ft"�i���� �E���P������$�[ �����G�����P�^ ����x���O�Gu
�� ����������� �f������f�f�f�f�f��U��WVS�E���D�u�EVP�]��������}� tk��X�󋻀   ���H  �{u ��   �Ct�EċKx1҅ɉȋ���u��u��u�SRP�E�WP�Q���}� t����P��B��PR� ���E�B��@ ��t!�{ ��u�Cx��t���P�R�����tO�e��[^_]Ð�t& �C|���E���   �E��x tY�H=�ȉMĈCt��Cu�X���H�����    ��'    �E���B�P��RP� ���e��[^_]Ít& ��'    ���u���4 �E����E�    � �P�    ����t���j �u����ȃ��M��n����Y� �	�R� ���*��uB��P� ���p�N�Ft"�I����� �E���P������$�Y �����'�����P�> ����x���O�Gu
� ������������ �f������f�f�f�f�f�����D$ �$�t$��������f�f�f�f��U��WVS�E���4�uVP��������}� tq��X�󋻀   ���N  �{u ��   �Ct�E̋Kx1҅ɉȋ���u�u�u�u�SRP�E�WP�Q ��,�}� t����P��B��PR�c} ���E�B��@ ��t!�; ��u�Cx��t���P�R�����tO�e��[^_]Ð�t& �C|���E���   �EȀx tY�H=�ȉM̈Ct��Cu�X���B�����    ��'    �E���B�P��RP��| ���e��[^_]Ít& ��'    ���u��2 �Eȃ��E�    � �P�    ����t���j �u����ȃ��M��n����� �	�� ���*��uB��P�@ ���p�N�Ft"�	���� �E���P�����$�PW �����������P�� ����x���O�Gu
�e �����������T �f������f�f�f�f�f��U��WVS�E���4�uVP�������}� tk��X�󋻀   ���N  �{u ��   �Ct�E̋Kx1҅ɉȋ���u�u�SRP�E�WP�Q$���}� t����P��B��PR�I{ ���E�B��@ ��t!�! ��u�Cx��t���P�R�����tU�e��[^_]Ít& ��'    �C|���E���   �EȀx tY�H=�ȉM̈Ct��Cu�X���B�����    ��'    �E���B�P��RP�z ���e��[^_]Ít& ��'    ���u��0 �Eȃ��E�    � �P�    ����t���j �u����ȃ��M��n������ �	��� ���*��uB��P�   ���p�N�Ft"������  �E���P�x����$�0U �����������P��� ����x���O�Gu
�E  �����������4  �f������f�f�f�f�f���D$� H	���D$��i f�f�f�f�f�S���\$�C�H	P�i �\$ ��[�<���f�f�f�f�f�f�S���\$�s � � �C$��[�f�f�f�f�S���\$�s ��� ZY�s P�>� ��[�S���D$�\$���t���s P�� ���C$������[Ít& �C$���uٸ�����ᐋD$�@ �D$��� VS�   ���D$ �\$�t$�L$��������C����t1҃�����RQ�v �l� ����u���v �� ������C����[^� f�f�f����D$�p �t$j�t$ �r� ���f��VS���\$�t$�s �t$jV�� ����~�T��S$��[^����������������C$������[^�f�����D$�T$���t �R �D$�T$���"� ��    ��'    ���r ��� �����������f�f�f��VS���t$�\$�T$��H�D$��@�uN��������C����jP�v �B� ����t����[^� f����v ��� ������C����[^� ���t$,j RPVS�у��؃�[^� f�f����D$� �p�P�t$�
������f�f�f�VS���t$��@�\|��tX�{ t$�C'��P�t$V�2  ��[^Í�    ��    ��S�, ����P�
   ����t�j
S�҃�����-� f�f�f�f�f�f��S���\$�C�H	�C    �C    �C    �C    �C    �C    P�� �D$$���C$�����C ��[�f�f�f��D$�@ �f�f�f�f�U��WVS�E��0�u�]�F    jVP�  ���}� �  �É߉E̋�@�\x�C;C�]��   � ���V���}ȍv ;E̍J�M���������������  �M�;M�  �]ԋ{�])ӍK��]ԋS)�9�Nу����   ����Q�u�W��� ��)���D�RW���u�� �}ԉ؉�]V��G;G�G�V�  � �_�����P��� ����X��K�C��  �I� �}��    1ҍ�&    ��'    �M��~�E�  �F��u,������x��WRW�t ���e��[^_]Ð��&    ��uӍe��[^_]�f����t+9E̺   u��EЋ}ԉF�G;G��   ��0҉G�f��   �v�����    �Mԋ]�}��A�Q���F9�sD���A9�sz� �V�}�\�����    ��    �}ԃ��W�P$���V�9�������'    �]ԃ��S�P(�����uS�V�}�����]ԃ��S�P$���������    ��'    �]ԃ��S�P$���Ë}ԃ��W�P(��1������]ԋC�S�M������S�����P�9� ���p�N�Ft�����}�҉��� ��S�MN �����������������x� ��S�/N f�f�f�f�f�f�f��U��WVS��,�}���  �E���@    jP�E�P� �E������   �}� ��   �E�}�]� �@�Dx�ǉEЋ@;G��  � �}���E� �uȋ��t& 9E�������ts9}��   �EЋu�P�X)���)�9�O�����   ���U�V�u�S��� �����U�)م��E�E����X�E9ډx��   �9E�������u��}� t�}�G�����    ��'    �����   9E��   �E�e�[^_]Ív �}���u��}�E��G   ��   ��������������������E��9ډx�~   �EЃ��X9�s�}��������t& �}Ѓ��W�P$�}�����������u�u�(� ���e�[^_]ËE�@=���t	�}���G�}ЋG;Gsf���G�3����}Ѓ��W�P(�����uU�E�x������]����E�U��� P�B��PR�p ��������}Ѓ��W�P$�������}Ѓ��W�P(�֋EЋX�P������u&��P�\� �E�}��� x�O�Gt@������P�6� �E�}��� x�O�Gu�� �f������� ��S�DK �������������s� ��S�*K f�f�f�f�f�U��WVS�E��@j �uP� ���}� ��  �E�u�]����� p���v��Oփ���lPS�U��Y �$�w=  �Eĉ$��_ �E�u��� �@�Dx�ƉE̋@;F��  � �u��E�    ���uȍ�    �U�9U���   �����   �}ĉƋO�ɉM��h  �}������������A  �ŰE�+EЋz�R���U�)�9�O���  �4�Eԍ_���;  9���  �G�U��� ��  �Eԉ���t& ��'    ��� ��  ��9�u�)���VW�u��� �}�u��uЋG�;G�G��  �U�9U�� ���������   �E�}��u�  �E� �P��D    ҃����;��P�� �E�u��� p�N�F��  �w� �MЅ�u �E�   � �up��VRV��m ���E�e�[^_]Ð�t& �E�}�  �E� �P��D    �UЅ�uк   볉���'    9���   �}���t& �;1�1ɈEԃ���tY�   �� t�=   �  �b  �� �Y  ��@�@  ���M�W�{e �M�����������'    ��Eԃ�u��EԄ���   �}���    ���m�������'    �E�E��ǍX���ü�F�V9��  ���F9��&  � �]�v�����    1����t& ��'    ����������   �� t�=   ��   w<�� �  ��@��   ���M�W�d �����M���	����������������=   ��   =  u~���M�W�)d �����M���	��p�����9�������}��q�����    ��'    =   ��   =  ��   ���M�W��c �����M���������&    ��'    1�	�������&    ���M�W�{c �����M���	������f����M�W��c �����M���	������f����M�W��c �����M���	�����f����M�W�c �����M��������t& ���M�W�{c �����M���������t& 1����������'    ���M�W�c �����M��������t& �ũ��V�P$���|����ũ��V�P(�����u8�]������[����ũ��V�P$���]�D����ũ��V�P$�������űF�V�����E�    ���1�����P�I� �E�u��� p�N�Ft�������� ��S�\E �����뺃��Ɖ�S�XZ ���������������s� ��S�*E f�f�f�f�f�U��WVS�E��@j �uP� ���}� u;�E�   � ��    �}x��WRW�i ���v ��'    �E�e�[^_]ËEj � �p�j �u�� X�E�u�]�Z����?� p�V����Oʃ�lPS�M���R �$�-7  �Eĉ$�Y �E�u��� �@�Dx�ƉEȋ@;F��  � �E�    ��t& �}ĉƋO�ɉM��]  �}�������������   �UȋE�+EԋJ�z�ʉM�)�9�O��r  �4�EЍ_����   9��I  �G�U��� �8  �EЉ������ �#  ��9�u��)�VW�u�� �}ȃ�uԋG�;G�G�i  �U�9U�� �4������u�E�}� �P��D    �   �b���f��E�}� �P��D    �Uԅ��b����   �8������&    9���   �}���t& �;1�1ɈEЃ���tY�   �� t�=   ��  ��  �� ��  ��@��  ���M�W��_ �M�����������'    ��EЃ�u��EЄ��i  �}���    �����������'    �E� �P�Z;X�w�x���~��S�u�� �E��� �P���E� =F�}  �uȃE��F�V9��4  ���F9�������}ȃ��W�P$���}�9}���������������E�}��}� �P��D    ҃��������f�1����t& ��'    ����������   �� t�=   ��   w<�� �  ��@��   ���M�W�^ �����M���	����������������=   ��   =  u~���M�W�	^ �����M���	��p�����9������}��q�����    ��'    =   ��   =  ��   ���M�W�] �����M����.�����&    ��'    1�	�������&    ���M�W�[] �����M���	������f����M�W�] �����M���	������f����M�W��] �����M���	�����f����M�W��\ �����M��������t& ���M�W�[] �����M����t����t& 1��i�������'    ���M�W�f] �����M����D����uȃ��V�P(�����uW�}�9}�������`������������������@�    �X�� �p����uȃ��V�P$������I����E�    �����}ȋG�W�Y�����uc��P�-� �E�u��� p�N�Ft=��������Ɖ�S�ST �������E�    ��E�    ������a� ��S�? ������P��� �E�M��� H�I�Au�-� �Mԅ�����������x������� ��S��> f�f�f�f�U��WVS�E��0�]j�uP�V ���}� u-�   �E�}��� x�WRW�Pc ���E�e�[^_]�f��Ej � �p�j �u蜵 �Ë}�މEȋE��� �@�\x�C;C��  � ��1��щU��}��&    9E�tv�S�K����?)�)�9�N΃��M���   ���u��u�R�U��f� �UЉƃ�)օ�Du�VR�u��� �C����;C�C��   � �����?��   ���u����t 9EȺ   �  ��������������f����   ������琉ƋE� �P�J;H��M�w�H���~���u��u��� �E��� �P���E� =F��   �C�S��9�sY���C9��R����t& ��'    ���S�P$�������?�>������&    ����7����   �5�����    ��'    ���S�P(�������   ������������U��@�    �P�� �d������C;Cs0���C��������������    ��    ���S�P$���������S�P(����1���u=��P��� �E�}��� x�O�Gt�����Ӊ��K� ��S�< ������P�� �E�]��� X�K�Cu�� �Y����C�S������`�������� ��S�; �D$�f�f�f�f�f��D$�@�@�f�f��D$�@�@�f�f��D$�@�@,�f�f���T$�D$�R�R0�� f�f�f�f�f�f���T$�D$�R�R4�� f�f�f�f�f�f���D$�@�@�f�f��D$�@�@�f�f��D$�@�@,�f�f���T$�D$�R�R0�� f�f�f�f�f�f���T$�D$�R�R4�� f�f�f�f�f�f���D$� H	�!l ��D$� �	�k ��D$�@�@$�f�f��D$�@�@%�f�f��D$� H�� �1��f�f�f�f�f�f��1��f�f�f�f�f�f����f�f�f�f�f�f�f�S�T$1��\$9�s��
�����9�u�[�f�f�f�f�f�f�f���D$� �	�1H ��D$� �	�!H ��D$� ���H ��D$� ���H ��D$� ����G ��D$� �	��G ��D$� �	��G ��D$� (	��G ��D$� (	�G �S���D$�\$$P�D$,�@�pS�c� ��(��[� f�f�f�f�f�S���D$�\$$P�D$,�@�pS�3� ��(��[� f�f�f�f�f�S���D$�\$$P�D$,�@�pS�� ��(��[� f�f�f�f�f�S���D$�\$$P�D$,�@�p$S��� ��(��[� f�f�f�f�f�S���D$�\$$P�D$,�@�pS�� ��(��[� f�f�f�f�f�S���D$�\$$P�D$,�@�pS�s� ��(��[� f�f�f�f�f�S���D$�\$$P�D$,�@�pS�C� ��(��[� f�f�f�f�f�S���D$�\$$P�D$,�@�p$S�� ��(��[� f�f�f�f�f�S���D$�\$$P�D$,�@�pS��� ��(��[� f�f�f�f�f�S���D$�\$$P�D$,�@�pS�� ��(��[� f�f�f�f�f�S���D$�\$$P�D$,�@�pS�� ��(��[� f�f�f�f�f�S���\$�{C ��	tL�C��t��P��� ���C��t��P�� ���C��t��P�� ���C$��t��P�� ���\$��[�3E f��S���\$�{C ��	tL�C��t��P�\� ���C��t��P�I� ���C��t��P�6� ���C$��t��P�#� ���\$��[��D f��S���\$�{d ��	t9�C��t��P��� ���C��t��P��� ���C��t��P��� ���\$��[�fD f�f�f�S���\$S�����\$ ��[鵰��f�f��S���\$S�����\$ ��[镰��f�f��S���\$�H	S�Lg �\$ ��[�o���f�f�f�f�f�f�f��S���\$��	S�f �\$ ��[�?���f�f�f�f�f�f�f��S���\$��	S�C �\$ ��[����f�f�f�f�f�f�f��S���\$��	S�|C �\$ ��[�߯��f�f�f�f�f�f�f��S���\$S�����\$ ��[鵯��f�f��S���\$�H�S� �\$ ��[鏯��f�f�f�f�f�f�f��S���\$���S��B �\$ ��[�_���f�f�f�f�f�f�f��S���\$���S��B �\$ ��[�/���f�f�f�f�f�f�f��S���\$S�����\$ ��[����f�f��S���\$��	S�|B �\$ ��[�߮��f�f�f�f�f�f�f��S���\$��	S�LB �\$ ��[鯮��f�f�f�f�f�f�f��S���\$�(	S�B �\$ ��[����f�f�f�f�f�f�f��S���\$�(	S��A �\$ ��[�O���f�f�f�f�f�f�f��S���\$�D$��)�RP�t$(�� ����[�f�f�f�f�f�f�f�U��VS�]���C�� 	P�f: �]���e�[^]�uA �ƃ�S�jA �4$�23 f�S���\$S�����\$ ��[鵭��f�f���D$� �	�����S���\$��	S�|����\$ ��[����f�f�f�f�f�f�f��U��VS�]���C���P��9 �]���e�[^]��@ �ƃ�S��@ �4$�2 f�U��VS�]�s� 	�
F 9�t��t��V��� ���C��t���P�R���C��P�W9 �]���e�[^]�f@ �ƃ�S�[@ �4$�#2 f��S���\$S�����\$ ��[饬��f�f���D$� 	�_ �S���\$�	S�|_ �\$ ��[�o���f�f�f�f�f�f�f��S���H�Y��ɉX~��[Ív ��'    ��RP�� ����[�f�f�f�f�f�f�f�U��WVS�E��,�}j P�u�u賿 �ÉE̍E��j P�u�u蚿 �K�P�ƉEȃ���UԉM�f���VSW�e� ����u^��S�	� �4$���� ���;]���;u�u+1ۄ��ËEȃ�=�Eu6�Ẽ�=�Eu>�e��[^_]Ä�uL����딍t& �ËEȃ�=�EtʍU�������Ẽ�=�EtU�������e��[^_]Ív ��'    �����녉ËẼ�=�Et�U�������S�Y0 f�f�f�f��VS�ƉӃ�P�! ����@=��u����[^Ív ��'    ��SV�Ѓ���[^�U��VS�]���C���P�7 �]���e�[^]�> �ƃ�S�
> �4$��/ f�U��VS�]���C���P��6 �$��= �]���e�[^]�=����ƃ�S��= �4$�/ f�f�f�f�f�U��VS�]���C���P�v6 �$�= �]���e�[^]�����ƃ�S�r= �4$�:/ f�f�f�f�f�U��WVS�E��,�]�}�u�Fj PVW�[� �P�)��E�6�ỦEԉ$蠳���uȉǃ����&    �u�VW�u�3� ��9E�w-����W�E��<� _�u��c������uԉ�VP�u�� ����PWS裴 �4$�� ���;u�ta����P�J;H��M�w�H���~���u�S�� ����P�� �=F�b����U��@�    �P�� �L�����    ��    ��W�� �Eȃ���=�Eu�e��[^_]� �U��3����e��[^_]� ����7�� �Eȃ�=�Et�U��������=�Et�U��������V�- ��P�a� �<$�� ���1������믉�릃�P�>� ����f�f�f�f��WV�z	S��j j�K �   �Ɖ��������8�u$�D$ ��P�t$$�t$ ��� ���É�[^_Ít& ��S�� �p�4$輱������VSP�)� XZhz	j� K �D$0��P�t$$�t$ �� Y^Wj����J �<$�H� ����[^_�f�f�f�f�f�f�f��UWVS���\$ �|$$�t$(�l$,�S��t��t,��@=��u8����)�PWU�� ����[^_]Í�&    ��S�7 ����@=��tȉl$,�t$(�|$$�\$ ��[^_]��f�f�f�f�f�f�f��UWVS���T$0�\$4�D$8�R��t��������[^_]Ð�t& ��1�1��FЉD$f��   �����tC����  wX����  ��   ����   ���G  ��V�H ������	ōt& ����u�����[^_]Í�&    ��'    ��   �  wb�� ��   ��@��   ��V�NH ������	�뫍t& ��'    ����   ����   ��V�MG ������	��v�����    ��   tH��  ��   ��V�G ������	��D����t& ��V�aH ������	��(������&    ��V��G ������	��������&    �|$	��	���������V��G ������	���������&    1�	��������&    ��V��F ������	��������&    ��V�F ������	��������&    ��V��G ������	��h���f�f�f�f�U1���VS�U�]���h 	�C    �����Cj j S�Y ���e�[^]Éƃ�S��7 �4$�) f�f�U1���VS�U�]���h 	�����C�E�Cj j S�BY ���e�[^]Éƃ�S�7 �4$�U) f�f��U1���VS�U�]���h 	�C    �����C�u�uS��X ���e�[^]Éƃ�S�:7 �4$�) f��D$��R����u�@�@Í�&    ��f�f�f�f�f�f�f��D$��R����u�@�@Í�&    ��f�f�f�f�f�f�f�S���D$$�\$ ��R����u'���T$R�@�pS�s� ���؃�[� ��&    ��PS�҃��؃�[� f�f�f�f�f�f��S���D$$�\$ ��R����u'���T$R�@�pS�� ���؃�[� ��&    ��PS�҃��؃�[� f�f�f�f�f�f��S���D$$�\$ ��R�� �u'���T$R�@�pS賺 ���؃�[� ��&    ��PS�҃��؃�[� f�f�f�f�f�f��S���D$$�\$ ��R��P�u'���T$R�@�p$S�S� ���؃�[� ��&    ��PS�҃��؃�[� f�f�f�f�f�f���D$��R ����u�@�@,Ð��&    ��f�f�f�f�f�f�f����T$$�D$ �
�I$����u�R�R0���� �v ��'    ��RP�D$�у��D$��� f�f�f�f����T$$�D$ �
�I(����u�R�R4���� �v ��'    ��RP�D$�у��D$��� f�f�f�f�U1���VS�U�]���( 	�C    �����Cj j S��T ���e�[^]Éƃ�S�<4 �4$�& f�f�U1���VS�U�]���( 	�����C�E�Cj j S�rT ���e�[^]Éƃ�S��3 �4$�% f�f��U1���VS�U�]���( 	�C    �����C�u�uS�T ���e�[^]Éƃ�S�3 �4$�b% f��D$��R���u�@�@Í�&    ��f�f�f�f�f�f�f��D$��R�� �u�@�@Í�&    ��f�f�f�f�f�f�f�S���D$$�\$ ��R����u'���T$R�@�pS�ӷ ���؃�[� ��&    ��PS�҃��؃�[� f�f�f�f�f�f��S���D$$�\$ ��R����u'���T$R�@�pS�s� ���؃�[� ��&    ��PS�҃��؃�[� f�f�f�f�f�f��S���D$$�\$ ��R����u'���T$R�@�pS�� ���؃�[� ��&    ��PS�҃��؃�[� f�f�f�f�f�f��S���D$$�\$ ��R���u'���T$R�@�p$S賶 ���؃�[� ��&    ��PS�҃��؃�[� f�f�f�f�f�f���D$��R ��0�u�@�@,Ð��&    ��f�f�f�f�f�f�f����T$$�D$ �
�I$��@�u�R�R0���� �v ��'    ��RP�D$�у��D$��� f�f�f�f����T$$�D$ �
�I(��`�u�R�R4���� �v ��'    ��RP�D$�у��D$��� f�f�f�f��L$�D$1҅�� �	�@    ���@    �@ �P�@ �@ �@    �@    �@    �@     �@$    �@(    �@,    �@0 �@1 �@2 �@3 �@4 �@5 �@6 �@7 �@C �f�f�f�f��L$�D$1҅�� �	�@    ���@    �@ �P�@ �@ �@    �@    �@    �@     �@$    �@(    �@,    �@0 �@1 �@2 �@3 �@4 �@5 �@6 �@7 �@C �f�f�f�f�U1���WVS�� �U�]���h 	�C    ���Cj j S�0Q �u�H	�z	�   ���t�u�@��   �u�e�[^_]Í�    ��'    �u��j �uV��' ��j �u�S��P �4$�	( ���e�[^_]É�������S�MR �4$��  ��S��. �4$��  f�f�U1���WVS�� �U�]���( 	�C    ���Cj j S�0O �u��	�z	�   ���t�u�@��   �u�e�[^_]Í�    ��'    �u��j �uV�' ��j �u�S��N �4$�9' ���e�[^_]É�������S�Q �4$�  ��S�,. �4$�� f�f��L$�D$1҅�� �	�P�f�f�f��S���D$�\$��t$<�t$<�t$<�L$<Q�t$<�t$<�t$<�t$<PS�R��4��[� f�S���D$�\$��t$<�t$<�t$<�L$<Q�t$<�t$<�t$<�t$<PS�R��4��[� f��L$�D$1҅�� �	�P�f�f�f��S���D$�\$��t$<�t$<�t$<�L$<Q�t$<�L$<Q�t$<�t$<PS�R��4��[� S���D$�\$��t$,�L$,Q�t$,�L$,Q�t$,�t$,PS�R��$��[� f�f�f�f�U1���VS�U�]�����C    �����Cj S�� ���e�[^]Éƃ�S�, �4$�f f�f�f�U1���VS�U�]���������C�E�Cj S�D� ���e�[^]Éƃ�S�O, �4$� f�f�f��U1���VS�U�]�����C    �����C�uS��� ���e�[^]Éƃ�S��+ �4$�� f�f���D$��R����u�@�@$Í�&    ��f�f�f�f�f�f�f��D$��R����u�@�@%Í�&    ��f�f�f�f�f�f�f�S���D$$�\$ ��R��@�u'���T$R�@�pS�3� ���؃�[� ��&    ��PS�҃��؃�[� f�f�f�f�f�f��S���D$$�\$ ��R��p�u'���T$R�@�pS�ӯ ���؃�[� ��&    ��PS�҃��؃�[� f�f�f�f�f�f��S���D$$�\$ ��R����u'���T$R�@�pS�s� ���؃�[� ��&    ��PS�҃��؃�[� f�f�f�f�f�f���L$�D$1҅�� �	�@    ���@    �@ �P�@    �@    �@    �@     �@$ �@% �@d �f�f�f�f�f�f��U1���WVS��$�M�]�����C    ���Cj S��� �u�H��z	�   ���t�u�@��   �u�e�[^_]����������������u��j �uV�/" XZ�u�S�d� �4$�\" ���e�[^_]É�������S�@� �4$�( ��S�O) �4$� f�f�f���L$�D$1҅�� ���P�f�f�f��S���D$ �\$��t$<�t$<�t$<�t$<�t$<�t$<�t$<PS�R��4��[� f�f�f�f�S���D$ �\$��t$<�t$<�t$<�t$<�t$<�t$<�t$<PS�R$��4��[� f�f�f�f�S���D$ �\$��t$<�t$<�t$<�t$<�t$<�t$<�t$<PS�R(��4��[� f�f�f�f�S���D$ �\$��t$<�t$<�t$<�t$<�t$<�t$<�t$<PS�R,��4��[� f�f�f�f�S���D$ �\$��t$<�t$<�t$<�t$<�t$<�t$<�t$<PS�R0��4��[� f�f�f�f��L$�D$1҅�� ���P�f�f�f��S���L$,�D$�\$�Q�L$,Q�t$,�t$,�t$,PS�R��$��[� f�f�f�f�f�f�S���D$�\$��t$,�t$,�L$,Q�t$,�t$,�t$,PS�R��$��[� f�f�f�f�f�S���D$ �\$��t$<�t$<�t$<�L$<Q�t$<�t$<�t$<PS�R ��4��[� f�f�f�S���D$�\$��t$,�L$,Q�t$,�t$,�t$,PS�R$��$��[� f�f�f�f�f�f�f�U1���VS�U�]��� 	�C    ���C��+ ���Cj S�;  ���e�[^]Éƃ�S�v& �4$�> f�f�f�f�f�f�f�U1���VS�U�]��� 	���C�E�C�+ ���Cj S�� ���e�[^]Éƃ�S�& �4$�� f�f�f�f�f�f�f��U1���WVS���U�]�}��� 	�C    ���C�2+ ����PW�ǿ ����u�s���uS�` ���e�[^_]Ð�t& ��W�[� ���E�$�	������u�E�WP�s� �U���S벉����s� ��S�Z% �4$�" ��P��� �C��9�t��t��P�� ��蚜�����f�f�f��T$�D$�J�I��R�R�P�f�f�f��T$�D$�J�I��R�R�P�f�f�f��T$�D$�J�I��R�R�P�f�f�f���f�f�f�f�f�f�f��T$�D$�J�I ��R�R$�P�f�f�f��T$�D$�J�I,��J�I0�H�J�I4�H�J�I8�H�J�I<�H�J�I@�H�R�RD�P�f�f�f�f���T$�D$�J�IH��J�IL�H�J�IP�H�J�IT�H�J�IX�H�J�I\�H�R�R`�P�f�f�f�f���T$�D$�J�Id��J�Ih�H�J�Il�H�J�Ip�H�J�It�H�J�Ix�H�J�I|�H�J���   �H�J���   �H �J���   �H$�J���   �H(�R���   �P,�f�f�f�f�f�f���T$�D$�J���   ��J���   �H�J���   �H�J���   �H�J���   �H�J���   �H�J���   �H�J���   �H�J���   �H �J���   �H$�J���   �H(�R���   �P,�f�f�f�f��L$�D$1҅�� ���@    ���@    �@    �P�@    �@    �@    �@     �@$    �@(    �@,    �@0    �@4    �@8    �@<    �@@    �@D    �@H    �@L    �@P    �@T    �@X    �@\    �@`    �@d    �@h    �@l    �@p    �@t    �@x    �@|    ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ƀ�    �f�f��L$�D$1҅�� �	�P�f�f�f��S���L$<�D$ �\$�Q�L$<Q�t$<�L$<Q�t$<�t$<�t$<PS�R��4��[� f��L$�D$1҅�� 	�P�f�f�f���L$�D$1҅�� (	�P�f�f�f���D$��B��f�f��S���D$ �\$��t$<�t$<�t$<�t$<�t$<�t$<�t$<PS�R��4��[� f�f�f�f�S���D$ �\$��t$<�t$<�t$<�t$<�t$<�t$<�t$<PS�R��4��[� f�f�f�f�S���D$ �\$��t$<�t$<�t$<�t$<�t$<�t$<�t$<PS�R��4��[� f�f�f�f�S���D$ �\$��t$<�t$<�t$<�t$<�t$<�t$<�t$<PS�R��4��[� f�f�f�f�S���D$ �\$��t$<�t$<�t$<�t$<�t$<�t$<�t$<PS�R��4��[� f�f�f�f��L$�D$1҅�� h	�P�f�f�f��VS1����T$�\$���� 	���C�$ �C��[^Éƃ�S�� �4$� f�VS1����T$�\$���� 	���C��# �C��[^Éƃ�S� �4$�b f��D$��B��f�f���D$��B��f�f��S���D$�\$��t$,�t$,�t$,�t$,PS�R��$��[� f�f��D$��B��f�f���D$� �f�f�f�f���D$� F� f��U��WVS�z	���]�uS������u��	�   �������8�t�u�@��   �u�e�[^_]Ís��V� ��j �uV�F ���e�[^_]Éƃ�S������4$�X f�f�f�f�U��WVS�z	���]�uS�F= �u�	�   �������8�t�u�@��   �u�e�[^_]Ís��V� ��j �uV� ���e�[^_]Éƃ�S�p< �4$�� f�f�f�f�VS1����T$�\$��������C��! �C��[^Éƃ�S� �4$� f�S1����T$$�\$��������C�D$ P�z �C��[�f��D$��B��f�f��S���D$�\$��t$�t$PS�R����[� f�f�f�f�f�f��D$��B��f�f��U1���WVS���U�]��������C�<! �u�C�z	����   �t�u�@��   �u�e�[^_]É���'    �s��V� ��j �uV�V ���e�[^_]É�������S�����4$�b ��S� �4$�Q ���h�E�C( �T$ ���;B�Js$����tj h`	h�
	P��� ����t	���艡 �� f�f�UWVS��8�D$T�L$X�l$h�\$`�D$�D$\�L$��lP�������L$;l$`��   ���ÉD$��&    �] ��  �؄��Z  ��%�!  �}9|$`��   �U��  �Є��N  ��Ot	��E�p  �}9|$`��   �m��.  �����   ���|$�D$D���L$X�|$T� SR�t$l�t$$�t$l�t$l�t$l�t$l�|$DW�P�D$H�L$x�T$D��0�	ىT$t�T$4�L$x����,��9l$`�#����D$�t$@�L$L�T$L�D$H�D$H�V���,��[^_]� �v ��'    ��R �T$�|$������   ���A�����.  �5���f����E u��|$�W;W��   ��G�m�����    ��'    ��R ����uS��t���  ���������[ ����uS��t��  ��������1�1�������t& �Ӊ�1������t& �L$�Ã�j PV�҃��L$듍�    �L$�T$��j PV�Ӄ��L$�T$닍�&    ��'    �L$��j RV�D$ �Ѓ����L$����������������������L$�PQ�R4��������d���f�f�UWVS�
   ��8�D$\�t$T�|$X�D$$�D$`�D$ �D$t��lP�����D$ ���|$dt�|$d�   f��E�1��D$    ��    ����  ����  �D$���k  1�1��|$���   8�u@�D$9D$dt�|$��  �|$d��  ��d�D$X�(�D$@�0�x��,[^_]� �t& �D$;D$ds����  �����   ���ȋT$��
  ����   �B�<	w��L� �lJЉ���;D$`�n����9D$\�b����gfff������)څ���t�F;F��   ���F������D$�������    ��    �L$�A;A�   � �D$1������f��F;F��   �8�������    ��    �F;F�  �8�'�����    ��    �T$��R ����u?<*������T$��
  �������t& ���V�P(���D������������������L$����j*P�t$�҃��L$륍t& ���V�P$�������   �T$1����-����   �����v �D$l��=����t& �T$���L$$�Q�P$�D$$������T$������   �D$    ��������&    ���V�P$�������������   �����1������D$;D$d������������   �������������`���f�f�f�f�f�f�f��UWVS��8�l$d�t$T�|$X�\$\�ElP�����D$�D$,    ���L$QUjh'  j �L$,Q�t$l�t$lWV�t$lP�����t$4�|$8��,�D$��uV�L$�id�������ɋL$`HŉA����   ���t@��t1�1��|$T�tA8�u�D$\��D$@�0�x��,[^_]� �v �D$\�뺍�&    �F;Fsh�8볍v �C9Cs1�볍t& �L$���S�P$������L$u޸   ���������������1����y����   �b�����    ��    ���V�P$�����tω��8���f�f�f�f���h�E�  �T$ ���;B�Js$����tj h�	h�
	P�9� ����t	������ �� f�f���h�E�c  �T$ ���;B�Js$����tj hp�h�
	P�� ����t	���詙 �Ĺ f�f���h�E�  �T$ ���;B�Js$����tj h��h�
	P虸 ����t	����Y� �t� f�f�U��WVS��X�]�Cd�u�����Ƌ ���@=@���  �Eʃ�P�F�p�E�P荗 ���EЍH�P���E�MĉS��  ��R�����E��C���Eċ�@=@���  �E˃��}�P�F�pW�4� ��j �u��u�W��n �Eԃ��P���E�  �E��S�C1���t�E�� �Eă�<}���C��@=p���  �Ẽ�P�F�p�E�P�Ŗ ���E؋P��=�E�S��  ��R�R����E��C���Eċ�@=p��  �E̓��}�P�F�pW�p� ��j �u��u�W�n �E܃���=�E�K  �E��C��@=���E  �E΃�P�F�p�E�P�E��� ���E��P��=�E�S ��  ��R詇���E��C ���Eċ�@=����  �Eσ��}�P�F�pW�Ǖ ��j �u��u�W�fm �E����=�E��  �E��C��@=����  �F�@$�C$��@=����  �F�@%�C%���u�����E��@���{&�5lD<t����   �Eċ �@=����   ��C&�F�G�F�G�F�G�F�G�F�G�F�G�F�G�F �G �Eč{J�5pD�@<t����   �Eċ �@=����   ��CJ�F�G�F�G�F�G�F�G�F�G�Ff�G�e�[^_]Ít& ���u��e�  �Eă�� �@=���D����V$WRV�u��Ѓ��f�����    ��    ���u��%�  �Eă�� �@=���h����VWRV�u��Ѓ��e�[^_]É���'    �}��VW�Ѓ��:�����&    ��'    �M���V�M�Q�Ѓ�������t& ��'    ��V�Ѓ��W���f���V�Ѓ��-���f��UЃ�VR�Ѓ�������&    ��'    �}ԃ�VW�Ѓ��M�����&    ��'    �}܃�VW�Ѓ��������&    ��'    �U؃�VR�Ѓ��|�����&    ��'    �U��h����S �����U��X����q����v �U��H����S�U����U��8��������v �H��y��ɉx�������E��PR�Rv �������v ��'    �x��O����H��@����E��P�u�� v �S���&��������v��P�D� �������Eԃ�=�Et�U�������S�� ���E�    �E�    ���u��© �E�����t��P诩 ���E���t���P蜩 ��떃�P�Ω ���E�    �E�    뮉��� �Q���2�O��I�C���G�� ��S��� �E�    ��P腩 ���p����E��=�Et�U�����������������ǋE܃�=�Et�U���������f����h�E�s �T$ ���;B�Js$����tj h|�h�
	P��� ����t	���蹒 �Բ f�f���h�E�# �T$ ���;B�Js$����tj h�h�
	P話 ����t	����i� 脲 f�f���h�E�� �T$ ���;B�Js$����tj h �h�
	P�Y� ����t	����� �4� f�f�U��WVS��h�u�FC�u�����Ë ���@=��#  �C�@�F��@= ���  �C�@�F��B =0���  �C�@,�F,�B=����  �E���P�C�p�E�P�� ���EȋP��=�E�V�  ��R菁���E��F���E���@=���#  �E����}�P�C�pW譏 ��j �u��u�W�Lg �Ẽ���=�E��  �E��V�F1���t�E�� �E���<}���F��@=����  �E�P�C�p�E�P�?� ���EЋP��=�E�V��  ��R�̀���E��F���E���@=���   �EÃ��}�P�C�pW�� ��j �u��u�W�f �Eԃ���=�E��  �E��F��@=����  �Eă�P�C�p�E�P虎 ���E؋P��=�E�V ��  ��R�&����E��F ���E���@=���:  �EŃ��}�P�C�pW�D� ��j �u��u�W��e �E܃���=�E�?  �E��F��@=���  �Eƃ�P�C�p$�E�P�E���� ���E��P��=�E�V(��  ��R�}���E��F(���E���@=��Q  �Eǃ��}�P�C�p$W蛍 ��j �u��u�W�:e �E����=�E�v  �E��F$��@$=@���   �C�@0�F0��@(=`���   �C�@4�F4���u������E��@���~8�tD<t��t8�E�� �@=��uF��F8�C�G�Cf�G�C
�G
�e�[^_]Í�&    ���u���  �E���� �@=��t��SWRS�u��Ѓ��e�[^_]Í�    ��'    �U���SR�ЋE����J����t& ��'    �U���SR�ЋE��������t& ��'    �}��SW�Ѓ�������&    ��'    �M���S�M�Q�Ѓ��>����t& ��'    �}܃�SW�Ѓ��������&    ��'    �U؃�SR�Ѓ��X�����&    ��'    �}ԃ�SW�Ѓ��������&    ��'    �UЃ�SR�Ѓ��r�����&    ��'    �}̃�SW�Ѓ��������&    ��'    �Uȃ�SR�Ѓ��o�����&    ��'    ��S�Ћ���'�����S�Ѓ�� ���f���S�Ѓ������f��U��h����V������U��X����N����v �U��H����V(�*����U��8����}����v �U��(����V �a����U����������v �U������V������U�������+�����   �	�   ���m�E�    �E�    �E�    ��P�C� �����u���� �E�����t��P�� ���E���t��P�ϡ ���E���t��P輡 ����|���Eԃ�=�Et�U��_������E�    �E�    끉���c����E�    �l����3� ��S��� �����ŋẼ�=�Et�U�������S脡 ���E�    �E�    �E�    �'������������P�U� ���T������g����b��������p����E��=�Et�U����������������������!�E܃�=�Et�U��v������+����&����!����������������������h���f�f�f�f����h�E�� �T$ ���;B�Js$����tj h@�h�
	P�y� ����t	����9� �T� f�f�U��WVS��h�u�FC�u�����Ë ���@=���#  �C�@�F��@=����  �C�@�F��B =����  �C�@,�F,�B=����  �E���P�C�p�E�P�"� ���EȋP��=�E�V�  ��R�y���E��F���E���@=���#  �E����}�P�C�pW�͇ ��j �u��u�W�l_ �Ẽ���=�E��  �E��V�F1���t�E�� �E���<}���F��@=����  �E�P�C�p�E�P�_� ���EЋP��=�E�V��  ��R��x���E��F���E���@=���   �EÃ��}�P�C�pW�
� ��j �u��u�W�^ �Eԃ���=�E��  �E��F��@= ���  �Eă�P�C�p�E�P蹆 ���E؋P��=�E�V ��  ��R�Fx���E��F ���E���@= ��:  �EŃ��}�P�C�pW�d� ��j �u��u�W�^ �E܃���=�E�?  �E��F��@=P���  �Eƃ�P�C�p$�E�P�E��� ���E��P��=�E�V(��  ��R�w���E��F(���E���@=P��Q  �Eǃ��}�P�C�p$W軅 ��j �u��u�W�Z] �E����=�E�v  �E��F$��@$=����   �C�@0�F0��@(=����   �C�@4�F4���u�����E��@���~8�tD<t��t8�E�� �@=��uF��F8�C�G�Cf�G�C
�G
�e�[^_]Í�&    ���u����  �E���� �@=��t��SWRS�u��Ѓ��e�[^_]Í�    ��'    �U���SR�ЋE����J����t& ��'    �U���SR�ЋE��������t& ��'    �}��SW�Ѓ�������&    ��'    �M���S�M�Q�Ѓ��>����t& ��'    �}܃�SW�Ѓ��������&    ��'    �U؃�SR�Ѓ��X�����&    ��'    �}ԃ�SW�Ѓ��������&    ��'    �UЃ�SR�Ѓ��r�����&    ��'    �}̃�SW�Ѓ��������&    ��'    �Uȃ�SR�Ѓ��o�����&    ��'    ��S�Ћ���'�����S�Ѓ�� ���f���S�Ѓ������f��U�舾���V������U��x����N����v �U��h����V(�*����U��X����}����v �U��H����V �a����U��8��������v �U��(����V������U������+�����   �	�   ���m�E�    �E�    �E�    ��P�c� �����u��� �E�����t��P�� ���E���t��P�� ���E���t��P�ܙ ����t���Eԃ�=�Et�U��������E�    �E�    끉���c����E�    �l����S� ��S�
� �����ŋẼ�=�Et�U��-�����S褙 ���E�    �E�    �E�    �'������������P�u� ���T������g����b��������p����E��=�Et�U�迼�������������������!�E܃�=�Et�U�薼�����+����&����!����������������������h���f�f�f�f����h�E�	 �T$ ���;B�Js$����tj h<�h�
	P虡 ����t	����Y� �t� f�f���h�E�� �T$ ���;B�Js$����tj h��h�
	P�I� ����t	����	� �$� f�f���h�E�s �T$ ���;B�Js$����tj h��h�
	P��� ����t	���蹁 �ԡ f�f�U��WVS��   �E�]�}(��L����E$��P����E��lP��T���������X��T����l������~ ����   �VB����d�������   ��ƅg��� ��e�����P�����f�����d�����h������u Ph�   ��WQ��� �����������!�%����t�������  DVD�L��� ����� )��҈�T���u%���VWS�P0��T�����9Ƹ   EȈ�T����E�����T����A�e��[^_]� ��&    ��P���ƅf��� ��e����:�����&    ����T���V��  ����%   ��T����@=���������j%V�Ѓ���T��������f�f�f�f�f����h�E� �T$ ���;B�Js$����tj h��h�
	P�	� ����t	����� �� f�f���h�E�3 �T$ ���;B�Js$����tj h`�h�
	P蹞 ����t	����y 蔟 f�f���h�E�� �T$ ���;B�Js$����tj h��h�
	P�i� ����t	����) �D� f�f�S��h�E� ���D$ ���1�;J�Zs!����tj h`	h�
	R�� ��������[�f�f�f��S��h�E�B ���D$ ���1�;J�Zs!����tj h�	h�
	R�ĝ ��������[�f�f�f��S��h�E�� ���D$ ���1�;J�Zs!����tj hp�h�
	R�t� ��������[�f�f�f��S��h�E� ���D$ ���1�;J�Zs!����tj h��h�
	R�$� ��������[�f�f�f��S��h�E�R ���D$ ���1�;J�Zs!����tj h|�h�
	R�Ԝ ��������[�f�f�f��S��h�E� ���D$ ���1�;J�Zs!����tj h�h�
	R脜 ��������[�f�f�f��S��h�E� ���D$ ���1�;J�Zs!����tj h@�h�
	R�4� ��������[�f�f�f��S��h�E�b ���D$ ���1�;J�Zs!����tj h<�h�
	R�� ��������[�f�f�f��S��h�E� ���D$ ���1�;J�Zs!����tj h��h�
	R蔛 ��������[�f�f�f��S��h�E�� ���D$ ���1�;J�Zs!����tj h��h�
	R�D� ��������[�f�f�f��S��h�E�r ���D$ ���1�;J�Zs!����tj h��h�
	R��� ��������[�f�f�f��S��h�E�" ���D$ ���1�;J�Zs!����tj h`�h�
	R褚 ��������[�f�f�f��S��h�E�� ���D$ ���1�;J�Zs!����tj h��h�
	R�T� ��������[�f�f�f��UW1�VS���|$(�L$$�T$4�?�L$1ɉ���\$,���\$������������������+l$09�~/�o���<}w&)�;L$�1  �D$(����+l$0�<����9�ы|$(�݋D$ �9T$0�|$t0�t$0�Ǎt& ��'    ���F���9ֈG�u��+t$0�D$ ����L$������tP�v �L$�|$�h��?������   ��1����������&    �2�L0��9�u���D5 ���u��L$�����tU��&    �\$�x��\$(���~R������1ۃ���    ��'    ��L��9�u��ڍ�����u���[^_]Ív ��'    ��������녉��"���f�f�f�f�f�f��UWVS���\$0�L$$�D$,�l$4�T$8�t$<��tM������SR)��t$8QPU���������)��)�)�RSP踋 ������[^_]Í�    ��'    ������SR�t$8QPU������� )���[^_]�f�f�f�f��VS���\$4�D$0�t$,��RP�t$(�t$(�D$4PV����)����$[^�f�f�f�f�f��U��WVS��h�E�EȋE�ƉEЋE�E��E����EϋE��lP�E��|����$�E�E���  �ǋE���@l�@�4�����E��?  �E �8�E��@88�  �uԋF0�E���v�@ �u��w�EċE��7�H���   9���  �����u�  ���&    �����  ��9�u����r  �6���E�FP�E�P�f �Mԉ���A,)҉U���   ���AIډ]����   �؃��j P�E��p�E�j P�_ �؃� ��E��EԋH�X�M��H�E܉M��H���x�E܃�P�[ �E܃����u�W�u��u�SP������ËE܃� �P���x�E܃�P�m[ �E܃�)Ë@��)�9���  �E�j RSP�yY �Eԃ��@,��~7�]ԃ��CP�E�P��j �E������H  ����s,P�E�P�h ���E�U܋uċ@r�ǁ�   ���}���  1�ƍ}����6�E�FPW�ge �E���]�@9Ɖ��E��}���!��E��U��E���)��ƀ;w#��$�������'    �Eą���  ��t& �E��9�u΃}�v�Eă���P�E���PW�Ig ���E��P�9U���  �}� �m  �E���P�E�)�Pj j W�E] �E��� �}� u�uȋ]����SPV�R0��9ËE��k  ��=�E�P  �E܃�=�Et����������&    �E�}��@    �EψEЋE�8�}Љx�e�[^_]� ��&    )����K�����&    �Mԋq$�A4�u��w�E�A(���E�t��E����7�H�������9߉�s��Eԉ}��߉u��ӉE��v ��'    �1�1��PЉEԉU�����tp�   ��t�� �D  �^  =   �  �}  =   �B  =  �J  ���uԉM��� ���M�����	ƍ�    ��    ����u������^  �}��E���)��Eԉ��P����v ��'    �E�@�����Eԃ��p�pW�ae �����������&    �}� u$���u�W��g �܍�    ��    �}� ��������u�VW�if 뷍�&    �E܃�PW�c 롐�Eԋ@������t& �E܃��u�WP�] �Eԃ��@,�����Eԃ��@9P�E���P�E�P�f �E܃�VWP�d ������t& ����   ��tr��t1�	�������t& �}�	��	������f���@uރ��uԉM��T� �����M���	������t& ��'    ��9������E��u��}��Eԉ������f����uԉM��� �����M���	��P������uԉM��� �����M���	��0������uԉM��i� �����M���	��������uԉM��� �����M���	���������uԉM��� �����M���	�������U��i������&    ��jD�Ə ��XZ�C    ��	�C    �C    �C �C �C �C    �C    �C    �C     �C$    �C(    �C,    �C0 �C1 �C2 �C3 �C4 �C5 �C6 �C7 �CC �u�S�=����E��WS�pl�=�  ����E������E���P�E�)�PW��c ���E������E���� PW�1e �,����U�贪�������E�����������*�F�UPShF�hx���s �E���=�Et�U��t����E܃�=�Et�U��_�����S�� ��P�͆ ���a����P輆 ��$�P����+� ��S��� f�U��WVS��h�E�EȋE�ƉEЋE�E��E����EϋE��lP�E��\����$�E�E���  �ǋE���@l�@�4�����E��?  �E �8�E��@88�  �uԋF0�E���v�@ �u��w�EċE��7�H���   9���  �����u�  ���&    �����  ��9�u����r  �6���E�FP�E�P�^ �Mԉ���A,)҉U���   ���AIډ]����   �؃��j P�E��p�E�j P��V �؃� ��E��EԋH�X�M��H�E܉M��H���x�E܃�P�S �E܃����u�W�u��u�SP������ËE܃� �P���x�E܃�P�MS �E܃�)Ë@��)�9���  �E�j RSP�YQ �Eԃ��@,��~7�]ԃ��CP�E�P�b �E������H  ����s,P�E�P��_ ���E�U܋uċ@r�ǁ�   ���}���  1�ƍ}����6�E�FPW�G] �E���]�@9Ɖ��E��}���!��E��U��E���)��ƀ;w#��$�������'    �Eą���  ��t& �E��9�u΃}�v�Eă���P�E���PW�)_ ���E��P�9U���  �}� �m  �E���P�E�)�Pj j W�%U �E��� �}� u�uȋ]����SPV�R0��9ËE��k  ��=�E�P  �E܃�=�Et���ئ�����&    �E�}��@    �EψEЋE�8�}Љx�e�[^_]� ��&    )����K�����&    �Mԋq$�A4�u��w�E�A(���E�t��E����7�H�������9߉�s��Eԉ}��߉u��ӉE��v ��'    �1�1��PЉEԉU�����tp�   ��t�� �D  �^  =   �  �}  =   �B  =  �J  ���uԉM��`� ���M�����	ƍ�    ��    ����u������^  �}��E���)��Eԉ��P����v ��'    �E�@�����Eԃ��p�pW�A] �����������&    �}� u$���u�W�_ �܍�    ��    �}� ��������u�VW�I^ 뷍�&    �E܃�PW�c[ 롐�Eԋ@������t& �E܃��u�WP�U �Eԃ��@,�����Eԃ��@9P�E���P�E�P��] �E܃�VWP�\ ������t& ����   ��tr��t1�	�������t& �}�	��	������f���@uރ��uԉM��4� �����M���	������t& ��'    ��9������E��u��}��Eԉ������f����uԉM��� �����M���	��P������uԉM���� �����M���	��0������uԉM��I� �����M���	��������uԉM���� �����M���	���������uԉM��� �����M���	�������U��i������&    ��jD覇 ��XZ�C    ��	�C    �C    �C �C �C �C    �C    �C    �C     �C$    �C(    �C,    �C0 �C1 �C2 �C3 �C4 �C5 �C6 �C7 �CC �u�S������E��WS�pl��  ����E������E���P�E�)�PW��[ ���E������E���� PW�] �,����U�蔢�������E�����������*�F�UPShF�hx���k �E���=�Et�U��T����E܃�=�Et�U��?�����S��� ��P�~ ���Y����P�~ ��$�P���� ��S��� f�U��WVS�u���D�E�EЋE �E̋E��lPV���  �4$�C�����P  �ǍD$����ÉE����  �u,�u(�u$j hZ�j S�]�E�S�����M߃� �E�Qj PS�I �E���Eԋ@���x��S�?L �E���E��G<t����   ��@=����   ���u��u��u��z ���}� tL�Ẽ�SP�u�u�u�u�u������E���P���Eu~��V���  �E�e�[^_]� ���&    �Ẽ�SP�u�u�u�u�u����벐��W�W�  ����@=���^����MċU��u��RQW�Ѓ��Z�����    ��    �H��Y��ɉX��q����E߃�PR�H ���\����������E��=�Et�U��=�����V��  �$��� f�f�f�f�f�f�S���|$  �\$�D$�L$$�T$(u5�����t$0RQ�t$,�t$,PS��������؃�[� ��&    ��'    �����t$0RQ�t$,�t$,PS�u������؃�[� f�f�f�f��UWVS���D$4�L$0�\$D�|$@�t$8�l$<�D$�A)�%�   �� ��   1҃�tC�T$��W�D$PV��y �T$�t$@)�Չ\$H�l$D��,[^_]�x ��    ��'    ����lQ�������x ����   �E :AJt.8AHt)8AMu��~�E8��   ta�Qu8�tY1��o���f��Ј�   ���\�������������������SU�V�w �D$�|$H�\$@�D$D��,[^_]�Ex ��    �E ���   �F��E�F�������t& ��P�D$��  �L$���-   ��@=����   �E 8��[����y �%����+   �ȉL$聟�����E �L$8��1����y ������0   �ȉL$�U���8E ������������L$�y ������x   ���)������E8��+����L$�y ������X   ���������E������j-Q�L$�Ѓ��L$�5���f�f�f�f�f�f�VS���t$ �\$0�3V�t$4�t$4�D$,P�t$8�����3��$[^ÐUWVS�|$$ �l$�L$�t$t0������f��ȃ��������)����D�шu��)�[^_]ËD$ ��J��@t4�D$ ��% @  �������T��    ������������u�뷉덴&    �����������D�u��f�f�f�f�U��WVS��H�Eh�E�EԋE�E̋E�E���  �ƋE���@l�@���;���   �M�G&��0�t$�EЋI����ȉMȃ�J���E��Ã�@����!E �Uǅ��E ����8�FE �ڃ�SQ�u�P�FP������ )ƀ �ÉE�MȍF�U���   ���
  �u ���S  ����   �}�W9�~/�J���)̍M�t$��QP�E����VWRP�u�����]�� ���}�G    �}̉�����u�Mԃ��SPQ�R0��9ظ   E��E�}ԉ��8���A�e��[^_]� ��    �W'�����]��b�����    ��    �\ �UǉMȃ��)܍]�t$SP�����V�u�G%P�w�w�u�K����Uǃ� �]���MȄ�������������U ��������}�@��   ��@�U����������L
�]�H�W*��������&    ��'    �W&�����]�������    ��    ��jh�f~ ��X�EZ�G    ��	��l�G    �G    �G �G    �G    �G    �G     �G$ �G% �Gd PW������E��VW�pl��  �;�������W*�����]���������P�#v ��<$�P����P����P�
v ����v ��S�8� f�f�f�f�U��WVS��,�E�u�} �]�E��E�E܋F��E�uW�U؍E�������WRV�u�u�uP�����E�]����E��E܉]�]�E�E�U��E�S�e�[^_]� �t& ��h�E��  ���EЋFl���@���E̋ ���u  ������   �x�P �}Ћ~9���   )׉U̍G���)��E؍L$��W���PQ�M��@r �Eԃ��F    �M؋U�%�   �� ��   �}� �U�u5���WQS�P0��9ǋU��n  ����U�R�u�S�P0�U܃�9��E��E܋u�]�E�E�U��E�V�e�[^_]� ��    ��'    �x�P�}Ћ~9��5����}� �F    ���������U�R�u�S�P0�U܃�9��E������v ��'    �}� �t�������U�R�u�S�P0�U܃��M�9���   ���WQS�P0��9��E��:�����    ��    ��jh�v{ ��X�Fl�U�Y�B    ��	�B    �B    �B �B    �B    �B    �B     �B$ �B% �Bd PR��������u��u��vl��  �Ẽ�� �����E���������P�:s �uȋ�4$�P���N����P�s ����s ��S�L� f�f�f�f�f�f�S���\$�t$,�D$,P�t$,�t$,�t$,�t$,S�������$��[� f�f�f�f�f�f�f��VS���D$�\$�L$ �t$$��R�� Nu-���t$,VQ�t$,�t$,PS�������؃�[^� ���&    ���t$,VQ�t$,�t$,PS�҃��؃�[^� f�f�f�f�f�f�f�U��WVS��H�Eh�E�EԋE�E̋E�E��[�  �ǋE���@l�@�4������  �C&��0�L$�ƉE��E����Mȋx����J���E���@����!��U�P�AWV�u P�����Mȃ� �ƉE�)����{ ��   �}� ��   �E�@9�~1�P���)ԍU�\$��RQ���S�uP�E�P�u�����u�� �ًE�@    �Ē���u�}ԃ��VQW�P0��9�   E؋E�}ԉ8�X�e�[^_]� ��t& �D  �   1����U���)čD$RQ�����P�u�S%�E�R�s�s�u������� �}� �Eȋu���-�����   �!����E �������}�@��   1��� @  �}��������D�u�A�C*��������t& ��jh�x Z��Y�@    � �	�@    �@    �@ �@    �@    �@    �@     �@$ �@% �@d �E��lPS�~����E��WS�pl��  ���������C*�����u��M�������P��o ��$�P���J����P�o ����1p ��S��� f�f�f�f�S���\$�t$,�D$,P�t$,�t$,�t$,�t$,S�8�����$��[� f�f�f�f�f�f�f��UWVS���\$@�|$<�t$8�k��%����  �C�D$���t$L�L$LQSWV�t$LP������D$$�L$(�k�Ɖ�0�	ȉǋD$L�0�x�D$L��8[^_]� VS���D$�\$�L$ �t$$��R��`Qu-���t$,VQ�t$,�t$,PS�u������؃�[^� ���&    ���t$,VQ�t$,�t$,PS�҃��؃�[^� f�f�f�f�f�f�f�UWVS���|$D �D$4�T$8�t$<�D$�T$tX�\$0�v ��'    j j
���|$�l$UW�z� �T���j j
UW�%� �у��D$	��T$uċD$0��)�[^_]ËD$@��J��@tG�D$@�\$0% @  �������T��t$�|$������������t$�|$���	�u�럋\$0���������������T$�L$���Ѓ��D��Љ������׉T$	ǉD$u��W���f�f�f�f�f��U��WVS��X�E�U$h�E�EȋE�UԉE��E�E��E �E��_�  �ǋE���@l�@���3���  �F&��@�\$�E��E����@�Eă�J���E���@��!UϋU�����+EЋE�UԉыU���8M�v�EЋU��؃� ���Mσ�Q�u��u�RP�C(P� ����� )À~ �ǉE�C(��   �}� �   �Uԅ��T  �E�   ��   �u�N9�~/�Q���)ԍU�\$��RP�E����SVQP�u�F����}�� �؋u��M���A    ��u�uȃ��WPV�Q0��9��   E؋E�}ȉ8�X�e�[^_]� �t& ��'    �N'�����}��e�����    ��    �T? ���)ԍU�\$RP�����S�u�F%P�v�v�u������ �}� �}��� ����E�   �����MЋ]ԉ�	�������}�@��   1��E� @  �]��������L�}�H�N*��������    ��'    �N&�����}�������    ��    ��jh�r ��X�EZ�F    ��	��l�F    �F    �F �F    �F    �F    �F     �F$ �F% �Fd PV������E��WV�pl�>�  �3���p����N*�����}��	�������P�Sj ��4$�P���#E����P�:j ����j ��S�h� f�f�f�f�S���\$�t$,�t$,�D$,P�t$,�t$,�t$,�t$,S������$��[� f�f�f�f�f��UWVS���D$$�\$ �L$0�t$8�|$<�l$4��R���Vu#WVUQ�t$<�t$<PS�P������؃�[^_]� �WVUQ�t$<�t$<PS�҃��؃�[^_]� �U��WVS��X�E�U$h�E�EЋE�ỦEċE�E��E �E���  �ǋE���@l�@�4������  �E��@�s&�L$�u��@����M��Eԃ�J���E���@����!���P�A(�u�V�u��u�P�h����M��� �ƉE�)���(�{ ��   ������   �E�@9�~1�P���)ԍU�\$��RQ���S�uP�E�P�u�����u�� �ًE�@    �EĄ���u�}Ѓ��VQW�P0��9�   E؋E�}Љ8�X�e�[^_]� ��    �D  �   1����U���)čD$RQ�����P�u�S%�E�R�s�s�u������E��� �u�������,����E�   �����EȋỦ�	������}�@��   1��E� @  �}��������D�u�A�C*��������&    ��'    ��jh�&o ��X�EZ�C    ��	��l�C    �C    �C �C    �C    �C    �C     �C$ �C% �Cd PS获���E��WS�pl���  ���������C*�����u��<�������P��f ��$�P���A����P��f ����Ag ��S��� f�f�f�f�S���\$�t$,�t$,�D$,P�t$,�t$,�t$,�t$,S������$��[� f�f�f�f�f��UWVS���D$$�\$ �L$0�t$8�|$<�l$4��R��PZu#WVUQ�t$<�t$<PS��������؃�[^_]� �WVUQ�t$<�t$<PS�҃��؃�[^_]� �U��WVS��(�]h�E�*�  �ǋ���@�4����t�e�[^_]�����������������jD�fm ZY�@    � �	�@    �@    �@ �@ �@ �@    �@    �@    �@     �@$    �@(    �@,    �@0 �@1 �@2 �@3 �@4 �@5 �@6 �@7 �@C SP�E��޼����W�u��3���  ����e�[^_]�����P�e ����?����P��d �U��$�P����ae ��S�� f�f�f�f�U��WVS��(�]h�E���  �ǋ���@�4����t�e�[^_]�����������������jD�6l ZY�@    � �	�@    �@    �@ �@ �@ �@    �@    �@    �@     �@$    �@(    �@,    �@0 �@1 �@2 �@3 �@4 �@5 �@6 �@7 �@C SP�E�������W�u��3��  ����e�[^_]�����P��c ���>����P��c �U��$�P����1d ��S�� f�f�f�f�U��WVS��(�]h�E���  �ǋ���@�4����t�e�[^_]�����������������jh�k ZY�@    � �	�@    �@    �@ �@    �@    �@    �@     �@$ �@% �@d SP�E��s�����W�u��3��  ����e�[^_]�����P��b ���=����P��b �U��$�P����6c ��S�� f�f�f�f�f�f��U��WVS�   ��T�E�}�E$�u �E��E�Wl�]�R�U��E��E�E��E�P������EċG���M؅��M�I؉���VQ��8  W��  ���G�CEƃ����)����  �t$�M��EԍEԃ��u�����u�SQj VP�ω���U����E�R�����]Ѓ��K���)̍L$����M��M��H����  ����  ��R������  ��SV�u��^ �]Ѓ��ڃ��U�Sj.V�H] �����U���   �M�)�E��I$��MĀy ��   �G9�~2�P���)ԍUЍ\$��R�u����SWP�E�P�u�R����UЃ� �]��E��G    ����u#�}����UċR�u�W�P0�Uă�9¸   E؋E�}��8�X�e�[^_]� ��EĀx �q�����~$�F<9�`����N��0��	�P���</�H���1��T���)ԍT$����U����+���   ��   1�1ۍUЋu�R�U��M�RQP�F%P�v�v�u����]Ѓ� �ډ]�������v ��'    ���E�P�T�  �E�����R�����n�����u�SVP�ҋ]Ѓ����l�����    �u����   �]л   ��u���a������]�SV�u��:\ ���U��+���f�f��S���\$�t$8�t$8j �D$<P�t$<�t$<�t$<�t$<S�������4��[� f�f�f�f��U��WVS�   ��T�E�}�u �E��E�WlR�U��E��E�E��E�P�����EċG���M؅��M�I؉���VQ��H  W�s�  ���G�C$Eƃ����)���  �t$�M��EԍE��u,�u(����u$SQj VP赆���U����E�R�Ʀ���]Ѓ��K���)̍L$����M��M��H����  ����  ��R������  ��SV�u���Z �]Ѓ��ڃ��U�Sj.V�.Z �����U���   �M�)�E��I$��MĀy ��   �G9�~2�P���)ԍUЍ\$��R�u����SWP�E�P�u�8����UЃ� �]��E��G    ����u#�}����UċR�u�W�P0�Uă�9¸   E؋E�}��8�X�e�[^_]� ��&    �EĀx �k�����~$�F<9�Z����N��0��	�J���</�B���1��T���)ԍT$����U����+���   ��   1�1ۍUЋu�R�U��M�RQP�F%P�v�v�u����]Ѓ� �ډ]�������v ��'    ���E�P�4�  �E�����R�����h�����u�SVP�ҋ]Ѓ����f�����    �u����   �]л   ��u���a������]�SV�u��Y ���U��%���f�f��S���\$�t$8�t$8�t$8jL�D$<P�t$<�t$<�t$<�t$<S�������4��[� f�f��S���\$���tN�C���t
��[Ð�t& �B;Bs� �C��[Í�    ��'    ���R�P$�����u��    ��[ø�����f�f�f�f�f�f��VS���t$ �\$$�����   1҃~�t!�����   1Ƀ{�t/8�����[^Ít& �P;Ps8��F1��͍�&    ��'    �H;Hs8�1ɉC8�����[^Ð�t& ���P�R$�����u��    �   �f��T$���P�Q$������T$u��   �    8�����[^ú   �E����   �M���f�f�f�f�f�f�U��WVS��(�E,��lP�ۢ���ǋE(����   ���)čE�\$��P�E���P���������t)����'    �E0��}�E�U����W�e�[^_]� �E��P�$������E(����t�1��]�1��M�U$���'��&    ����U�PW�Q��8E�U�t��;u(t��� :E�uՋE܉4�����;u(u�؉]��E�    ���]��  ��    ��    ��}$���   �4��X �ǉ؃����ǋ��U$���4��X ��9�G؃�;u�r߉��߉ËE��t�P;P�\  ���P�E�����E��E�9�������E��P�EP�������������1��u�����    8E�tK����9։vF�<��M$����M���M�ɈE���   �E���uǋA;A��   � 8E�Eu���9�w����u�������}��C����E��t��P���  �E��������}$���u��<��E���W��V ��9���v��    �E��P�EP��������t`9�������E �}��8������t& ����U�Q�P$������U��M����E    �����������������������P�R(�������7�M��Q�E��������8E�u��E��t��P���  �E��������9��I����[���f�f�U��WVS�]��8�E,��lP�ȟ���E܋E(����   ���)čD$������ǍEPS���������o  �]1��E�    �E�    ������������������  �E�����   �U��t-1�1��}��  8��  �U���  �E����8  �EӅ��  1��E�    �}�����������������E���9�vH�]���    �M$�<E܋�}؋��M�;sӋ}��M�8;tW�]����M؋}�9֋�����w�9uԋ}��}   �]��t�C;C��   ���C�E�����E��������&    ���o������&    �C;Cs� �U�E�����������f��B;B��   � �E1�8����������  ��t~�E0��}�E�U����W�e�[^_]� ��    �B;B��   � �E�������S�P$������o����E    �U��t��   �Y������S�P(�]�������E܋u�90t	9p�o������+U(9E(FU ��^������R�P$������(����E    �   �������R�P$������R����E    �E���������1�S1���������E(����E���   �}؉ʋ}$�,����'    �U��U܃��
PR�Q�U���8�t��;]�t��� 8�uӋE؉�����;]�u���}؋]��   ��t��S��  �]�E��������   1҉]��Ӄ��)čD$����E�E܍v ��'    ���U$���4��R �U������9�uߋ]��E�   ������E܋u�90���������E��������]�E�    �E�    �����E�    �E�    �{���f�f�f�f�f��UWVS��h��$�   �t$|��$�   �hlU莻���É,$贛���C�PH�T$(�PL�@P�T$,�D$0�C�@T�D$4�C�@X�D$8�C�@\�D$<�C�@`�D$@�C�@,�D$D�C�@0�D$H�C�@4�D$L�C�@8�D$P�C�@<�D$T�C�D$$    �@@�D$X�C�@D�D$\�D$���T$R��$�   j�T$(R�T$$R��$�   ��$�   ��$�   ��$�   ��$�   P������D$4�T$8��$�   ��$�   ��$�   ��$�   ��,�D$��uO�T$��$�   �P����   ���tD��t1�1���$�   �tB8�u
��$�   ���n��\[��^_]� �v ��$�   �볍t& �C;Csh�(믍v �G9Gs1�벍t& �T$���W�P$������T$u޸   ���������������1ۅ��x����   �^�����    ��    ���S�P$�����tω��4���f�f�f�f�UWVS��   ��$�   ��$�   ��$�   �hlU�h����É,$莙���C���   �T$0���   ���   �T$4�D$8�C���   �D$<�C���   �D$@�C���   �D$D�C���   �D$H�C���   �D$L�C���   �D$P�C���   �D$T�C���   �D$X�C���   �D$\�C�@d�D$`�C�@h�D$d�C�@l�D$h�C�@p�D$l�C�@t�D$p�C�@x�D$t�C�@|�D$x�C���   �D$|�C���   ��$�   �C���   ��$�   �C���   ��$�   �C�D$,    ���   ��$�   �D$���T$ R��$�   j�T$0R�T$,R��$�   ��$�   ��$�   ��$�   ��$�   P�5����D$4�T$8��$�   ��$�   ��$�   ��$�   ��,�D$��uV�T$��$�   �P����   ���tK��t1�1���$�   �tI8�u
��$�   ���n�Č   [��^_]� ��&    ��$�   �묍t& �C;Csh�(먍v �G9Gs1�뫍t& �T$���W�P$������T$u޸   ���������������1ۅ��q����   �W�����    ��    ���S�P$�����tω��-���f�f�f�f�UWVS��h��$�   �XlS詶���$��1��͖��Y��$�   ���M ���T$x�$�D$    ��    ��    ����   �|$|���  ��$�   ��t1�1Ƀ�$�   ���   8���   ;$�D$��   ����   ��$�   ������  ���d  ��%��   ��$�   �{�L��  �Ȅ���  ��O�D$    �Y  ��E�P  ����A��8�r  ���$������&    ���R�P$�������   �D$x    ��$�   ��t51Ƀ�$�   ��   �#����H;H�w
  �1ɉ�$�   8������D$��u;$t
��$�   ��t$p�D$x�T$|����V��\[^_]� ���������������T$x����g  �D$|�����   8���   �L$���_������������������B;B����� �D$|�K������&    �U �R �����.  ��t���  ���x�����    ��    ��$�   ���<��=  ����������U �R �����.
  ����   ��=  ���j������&    �B;Bsh�8���|$|8��+����B;B��	  ���B�D$|�����T$x�����t& �U �R �����.	  ��uZ�L$�T$x��������v ��'    �L$���R�P$������L$��	  �D$x    1Ҁ������������v ��'    ��  ������f��L$��j PU�҃��L$������&    ���o�������'    �F���p��&    ��$�   �D$(P��$�   ��$�   ��$�   ��$�   ��$�   ��$�   �D$4P� ����D$4��$�   �D$8��$�   ��,���������$�   P����������=  ���\  ��	t@�L$�T$x������&    ����$�   P�P���������=  ����  ��
u��T$x���r�����R�`�  Ǆ$�   ������$�   ���O�����    �D$P��$�   jjj�D$0P��$�   ��$�   ��$�   ��$�   ��$�   �D$4P�����D$4�T$8��$�   ��$�   ��,�D$��������D$��$�   �T$x���G�������    ��'    ����$�   P�`�������Pj U��r��������  ��$�   �x�D$x��t��P�k�  Ǆ$�   �������D$P��$�   jj	jW�(���&    �D$P��$�   jjj��$�   ��P�v ��$�   ��$�   ��$�   ��$�   ��$�   �D$4P�����������&    ��'    �F���p����f��F���   �T$ ���   �T$$���   �D$(�F���   �D$,�F���   �D$0�F���   �D$4�F���   �D$8�F���   �D$<�F���   �D$@�F���   �D$D�F���   �D$H�F���   �D$L���D$P��$�   j�D$0P��$�   ��P��$�   ��$�   ��$�   ��$�   ��$�   �D$4P�����������&    �F�PH�T$ �PL�T$$�@P�D$(�F�@T�D$,�F�@X�D$0�F�@\�D$4�F�@`�D$8���D$P��$�   j�D$0P��$�   ���a����t& ��'    ����$�   P� �������PjU�p��������������|$W��$�   jh�D�D$4P��$�   ��$�   ��$�   ��$�   ��$�   �D$4P�����D$4�T$8��$�   ��$�   ��$��$�   P��$�   P� �������������T$��������D$ �����������$�   P�]����D$���} ��  �EJ8D$t/����$�   P�2����D$���} ��  �EH8D$�F���W��$�   jjj �D$4P��$�   ��$�   ��$�   ��$�   ��$�   �D$4P�3����D$4�T$8��$�   ��$�   ��,W��$�   jj;j �|$4W��$�   ��$�   RP��$�   �D$4P�����D$4�T$8��$�   ��$�   ��,�������&    �F���p�R���f��|$ Whx�ho�U�+n��XZW�3����v �D$P��$�   jj=j ��$�   �2���f��|$ Who�hi�U��m��YXW������v �D$P��$�   jj;j ��$�   ��P�������&    ��'    �D$P��$�   jjj��$�   ��P������&    ��'    �D$P��$�   jjj ��$�   ��P������&    ��'    �|$ Whi�h`�U�;m��XZW�C����v �D$P��$�   jh'  j �D$0P��$�   ��$�   ��$�   ��$�   ��$�   �D$4P�Y����D$4�T$8��$�   ��$�   ��,�L$�������T$��$�   �Jd�������ҋT$xH��G��������������������F�Pd�T$ �Ph�T$$�@l�D$(�F�@p�D$,�F�@t�D$0�F�@x�D$4�F�@|�D$8�F���   �D$<�F���   �D$@�F���   �D$D�F���   �D$H�F���   � �����&    ��'    �F�P,�T$ �P0�T$$�@4�D$(�F�@8�D$,�F�@<�D$0�F�@@�D$4�F�@D�k������������������T$���P�Q$������T$�n���Ǆ$�       �   �m�����    ��'    �L$����j PU�҃��L$�����D$P��$�   jjj
��$�   ��P�b����U �J ����uz���������=  ������U �J ����uC���������=  �����v ��'    ����j PU�҃��������R�P(�����������j PU�у���몃���j PU�у����p����-   ����f���I����+   ����f���c���8��T$x�D$|����������������f��UWVS��(�l$T�t$D�|$H�\$L�ElP�`����@�L$���p�t$\�t$\U�t$\�t$\WV�t$\Q�v����t$4�|$8��,��������   ���t:��t1�1��|$D�t;8�u�D$L��D$0�(�H��[^_]� ��    ��'    �F;FsX�빍v �C9Cs1�빍t& �T$�$���S�P$������$�T$uظ   뎉���'    1��t��   �l����<$���V�P$������$tى��H���f�UWVS��(�l$T�t$D�|$H�\$L�ElP�@����@�L$���p�t$\�t$\U�t$\�t$\WV�t$\Q�V����t$4�|$8��,��������   ���t:��t1�1��|$D�t;8�u�D$L��D$0�(�H��[^_]� ��    ��'    �F;FsX�빍v �C9Cs1�빍t& �T$�$���S�P$������$�T$uظ   뎉���'    1��t��   �l����<$���V�P$������$tى��H���f�U��WVS��X�E �XlS�[����E�X�E�ZSP�\����H �p8���E��E� �u���t	�@(���E��E��E�F�x t�E܃�j P� ���E����E�Fj P�� �E��E�    ���E� �E�    �E�    �E� �p9�@4�u�1��E�EĀ|���   ��&    �D��$����t& �E��}���  �   �U����  �E����  �U���P  1�1��}���  8��  �}� ��  �Eă�����  �EċEĀ|��{����t& ��'    �E��ύv ��'    �U����   ��t& �E����D  �U��t-1�1��}���   8���   �U���D  �E����P  ������j
P�u��z9 �����R  +E��tD�<�E��P�Z;X�w�H���~�E���SP�s �E����P����E�=F�  ���U��t-�B;B�  ���B���E�����,�����    ��    �U��t91��}��   �)������&    �B;B�4  � �E1�8������t& �E��E��H���y�����&    ��'    �]�}�E$���WS����������B	  �E�u�U��E��V��=�E�q
  �E܃�=�E�K
  �E�e�[^_]� f��E̋x ���  �E̋@(���9  �E����E��������t& �E �@��  �}���  �Eą���  ����  �}��E�������E�<��  �}� t<��  �   �����v �E��P�EP����������  �}��E� �����}���"EЄ��^  �}� ������t& ��'    �E��x�v7�E���j j0P� ����t ���u	�E��@����P�E�j P�� ���}� t\�E��P�����  �E���P�	 �E����80t7�H���x�E���P�b	 ���E���j-jj j P�{ �E��� �@������E܋@��t:�}� �U������]�E�PS� �Ẽ�S�p�p蕝  �����]  �}� t�E̍]�}9p,������E���P�u(���  ���]�}������t& �B;B��  � �U�E��������v �U���s  �E���u�B;B�a  � �E�؋M��Q���:  ����������������U����  �U�������1��}��   �r����B;B�  � �E1��Y�����    �B;B��  � �U�E��������U�������������������������'    �B;B��  � �E��������'    �}�8_u(�}� u"�_,���W����u��E�1����������'    �Èx �3���8X�*����}� � ������E  �������E�VP�� ��1�������    ��    1�1ɈEԉ���'    ����tS���� t�=   ��   wS�� ��   ��@��   ���M�S�ܪ �M��������v ��'    ��Eԃ�u��Eԉ��\����v ��'    =   ty=  uB���M�S�M� �����M���빉���'    ���M�S�� �����M���뗍�&    1�댍�    ��    ���M�S薪 �����M����d����t& ���M�S�;� �����M����D����t& ���R�P$�����������E    �   �-����v ��'    ���R�P$����������E    �t������������������@�    �X�� �������    ��'    ���R�P(���U�������    ��    �B;B�1  ���B�E�����e���f����R�P$������:����E    ���������������������R�P$�����������E    �   �����v ��'    ���R�P$����������E    ���������������}� �	  �t& ��'    �E�1ۋ@�EԋEf�����   �}���   �E��t1�1҃}���   ��8���   ;]�������E��P�����}̃��W8��   ��� ����E �@�����E������v ��'    ���P�R$�����uZ�E    �E��t/1҃}��   �w����P;P��   ��E1҉�8��c���;]�u��H������&    �P;Ps���E������    ��'    �E��t�P;Ps!���P�E�������������    ��    ���P�R(���E�������������������P�R$������Z����E    �   �����v ��'    ���R�P$�����������E    ����������E��P�>�������Pj �u��]������������E���������P�N�  ���E�����E������E��P�EP�[���������   �E̋x(��u�E̋P ��������E��E�������E��P�EP���������W  �E̋X ��������E̋X(��t��������R�P(����������������������E� ������E��P�N����}̃��W8�]����E̋@ �E��E���Y�����P�`�  ���E�����E������E$������}�������}��� ���������}� �E���   �@$�EЍ]�}�E�   ��&    ��WS�&����U���9U���8�r�M�9M��0����e�����t& ��S�����MЋUԃ�8uӋU��t�B;Bs���B�E�����E�뗋��R�P(����E��P�=����}̃��W$8������E̋@(�E��E���P�����P�O�  ���E�����E��E�������@�E������E$������80�*����F����U��U���E�e�[^_]� �U��U����������ËE���=�Et�U��wU���E܃�=�Et�U��bU����S�� f�f�f�f��U��WVS��X�E �XlS�y���E�X�E�ZSP������H �p8���E��E� �u���t	�@(���E��E��E�F�x t�E܃�j P�^
 ���E����E�Fj P�F
 �E��E�    ���E� �E�    �E�    �E� �p9�@4�u�1��E�EĀ|���   ��&    �D��$����t& �E��}���  �   �U����  �E����  �U���P  1�1��}���  8��  �}� ��  �Eă�����  �EċEĀ|��{����t& ��'    �E��ύv ��'    �U����   ��t& �E����D  �U��t-1�1��}���   8���   �U���D  �E����P  ������j
P�u���+ �����R  +E��tD�<�E��P�Z;X�w�H���~�E���SP�� �E����P����E�=F�  ���U��t-�B;B�  ���B���E�����,�����    ��    �U��t91��}��   �)������&    �B;B�4  � �E1�8������t& �E��E��H���y�����&    ��'    �]�}�E$���WS���������B	  �E�u�U��E��V��=�E�q
  �E܃�=�E�K
  �E�e�[^_]� f��E̋x ���  �E̋@(���9  �E����E��������t& �E �@��  �}���  �Eą���  ����  �}��E�������E�<��  �}� t<��  �   �����v �E��P�EP�0��������  �}��E� �����}���"EЄ��^  �}� ������t& ��'    �E��x�v7�E���j j0P���  ����t ���u	�E��@����P�E�j P�3�  ���}� t\�E��P�����  �E���P���  �E����80t7�H���x�E���P��  ���E���j-jj j P���  �E��� �@������E܋@��t:�}� �U������]�E�PS� �Ẽ�S�p�p��  �����]  �}� t�E̍]�}9p,������E���P�u(�C�  ���]�}������t& �B;B��  � �U�E��������v �U���s  �E���u�B;B�a  � �E�؋M��Q���:  ����������������U����  �U�������1��}��   �r����B;B�  � �E1��Y�����    �B;B��  � �U�E��������U�������������������������'    �B;B��  � �E��������'    �}�8_u(�}� u"�_,���W����u��E�1����������'    �Èx �3���8X�*����}� � ������E  �������E�VP�6	 ��1�������    ��    1�1ɈEԉ���'    ����tS���� t�=   ��   wS�� ��   ��@��   ���M�S�,� �M��������v ��'    ��Eԃ�u��Eԉ��\����v ��'    =   ty=  uB���M�S蝜 �����M���빉���'    ���M�S�[� �����M���뗍�&    1�댍�    ��    ���M�S�� �����M����d����t& ���M�S苜 �����M����D����t& ���R�P$�����������E    �   �-����v ��'    ���R�P$����������E    �t������������������@�    �X�� �������    ��'    ���R�P(���U�������    ��    �B;B�1  ���B�E�����e���f����R�P$������:����E    ���������������������R�P$�����������E    �   �����v ��'    ���R�P$����������E    ���������������}� �	  �t& ��'    �E�1ۋ@�EԋEf�����   �}���   �E��t1�1҃}���   ��8���   ;]�������E��P������}̃��W8��   ��� ����E �@�����E������v ��'    ���P�R$�����uZ�E    �E��t/1҃}��   �w����P;P��   ��E1҉�8��c���;]�u��H������&    �P;Ps���E������    ��'    �E��t�P;Ps!���P�E�������������    ��    ���P�R(���E�������������������P�R$������Z����E    �   �����v ��'    ���R�P$�����������E    ����������E��P��������Pj �u���O������������E���������P螜  ���E�����E������E��P�EP����������   �E̋x(��u�E̋P ��������E��E�������E��P�EP�k��������W  �E̋X ��������E̋X(��t��������R�P(����������������������E� ������E��P�����}̃��W8�]����E̋@ �E��E���Y�����P谛  ���E�����E������E$������}�������}��� ���������}� �E���   �@$�EЍ]�}�E�   ��&    ��WS�v����U���9U���8�r�M�9M��0����e�����t& ��S������MЋUԃ�8uӋU��t�B;Bs���B�E�����E�뗋��R�P(����E��P�����}̃��W$8������E̋@(�E��E���P�����P蟚  ���E�����E��E�������@�E������E$������80�*����F����U���G���E�e�[^_]� �U���G����������ËE���=�Et�U���G���E܃�=�Et�U��G����S�iy f�f�f�f��U��WVS�UЃ�,�}  �u�}�E$�E�Ftn�M���Q�u(P�u�uWV�uR�b�����,�uЋ}��t�  �]�E�S�u(�u,�u��~ �E���0�x�E��P���Eu6�E�e�[^_]� ����'    �M���Q�u(P�u�uWV�uR�����f��p��~����x����SR��  ��뮉ËE���=�Et�U��F����S�tx f�f�U��WVS��8�E$�] ��lP�k�����ۉ��E�F�E�te�U��R�u(�u$�u�u�u�u�uP�c����EЋUԃ�,�E�E�U�X��uZ�}�M�P�]���E��_��   �E�e�[^_]� �U��R�u(�u$�u�u�u�u�uP����뙍�    ��    ��j S�u,��  �E,��� �ǋ@���x���u,��  �E,��� �ǋE�E��F<t��t*��@=��u^��S�u�W�{ �E���<�����    ��V�R  ����f��H��Y��ɉX��2����E��PR��  �������v ��'    W�}��SWV�Ѓ��E�������ËE��=�Et�U��E����S��v f�f�f�f�f�U��WVS1ۃ�4�E ��lP�E�P�Ž����X�EZP�EP�d��������E��F  �V�E�    1��E���t& ���E�F�  �Fd���E��  �}� ��  �E� �E� �C�<	��   ����S�u(���  ���   �E����  �P;P�'  ���E�����P�P;P�>  ��U�E����  1�1��}��[  8��o  �]�K��t-�Eԍ}��8E���  ��W�v�v�;�  ������  �E�}�U��C�W=�E�J	  �E�e�[^_]� ��&    8^$�G  8^\t8^bu���8M��{�����je�u(���  �E������  �P;P�  ���E�����P�P;P��  ��U�E��t1�1��}���   8��  �E��P�3�����8FK����   8FJ�E��x����-   ��P�u(�W�  �E���E����������t& �U�������1��}��   ������B;B��  � �E1�8�������E��P������������f��+   ������    �B;B��  � �E1��0�����&    �Eԃ�:E��������j.�u(��  ���E��������&    ���P�R(�E���E�������2����P;P�������    ���P�R$�����������E    ����������������������P�R$������l����E    �U����  �   �\������������������}� �w  �FN�E� �E� �E��F��t	:^%��   :^$�N  ����j
P�u��z ������  +Eȃ���0��P�u(��  �E����   �E����   �P;P�J  ���E�����P�P;P�a  ��U�E��t1�1��}���   8�������E��P��������F�����J���:^%�A����Eԃ�:E���  �EЅ��(  ����P�E�P���  �E���E� �E�    ���N����t& �U���>���1��}��]��o����B;B�	  � �E1��V�����    ��    �E$�    �2���f��Eԃ�:E��P  �E�@��t�EЃ�P�E�P�E�  ����j.�u(�5�  ���E���������'    :^\t	:^b�������:E�������}� u�E�X��t�EЃ�P�E�P���  ����je�u(���  �E����t�P;P��  ���P�E�����E��P�EP�ÿ��������  �E��P�<�����8FK����t8FJt�F�E�������    ��'    �V��t	8F%�  8F$�  ���������+P�u(�/�  ���E������v ���P�R(�E���E�������B����P;P�������    ���P�R$�����������E    ���������������������P�R(�E���E�����������������    ��'    ���R�P$�����������E    �E��5����t& ��'    ���R�P$������6����E    �   �����v ��'    ���E��Q�����t& �}ԉ��E�F�}ЉύE��j P��  �����������'    �E��P蔽������8^K����   8^J��   �V1�1��Mԉ���    ��'    ��t8F%t�8F$�.  �^N8��"  ����  �E�E�����  �P;P��  ���E�����P�P;P��  ��U�E���!  1�1��}���   8��  �E��V�   �E��E��������&    �]�C��������E���������&    �V��t	8^%�:  8^$�������������+P�u(��  �E����t��P蜎  �E�������E��P�EP貼�������Q����E��P�+����V�������]�S���!�����EЃ�P�E�P���M�  ���]������f��B;B��   � �E1�8�������E��P�Ȼ���V�   ���W�����&    ��j0�u(���  �E���E����f�����U��������   �����t& ��'    ���P�R(�E���E������tƋP;P�D����v ��'    ���P�R$������(����E    �f��}ԉÉ}Љ��A��������M�R�P$������M������E    �   ������v �E��W�����&    ���P�R(���U��������������������R�P$����������E    �   �C����U��b:���E�e�[^_]� �E(j � �p�j �u(�A�  ���E� �.����   ������ËE��=�Et�U��:����S��k f�f�f�f�f��U��WVS�u���4�E�F�]j V�R�  �EЉ4$�u$�u �u�u�u�u�uP������EЋUԃ�,�E�U��~  �u�E�V�u$�u(�u��n �E������   �}�tD��t1�1��}�tF��8�u�E$��}�E�U��E��W�P���Eu^�E�e�[^_]� ��P;Ps��E묋C9CsX1�뮍t& � ���u�P$�����u��E    ��t��   �z������&    �H��Y��ɉX����VR��  ��농t& ���S�P$�����u��   �?����ËE���=�Et�U��8����S�Uj f�f��U��WVS�u���4�E�F�]j V���  �EЉ4$�u$�u �u�u�u�u�uP�Q����EЋUԃ�,�E�U�]}  �u�E�V�u$�u(�u��hn �E������   �}�tD��t1�1��}�tF��8�u�E$��}�E�U��E��W�P���Eu^�E�e�[^_]� ��P;Ps��E묋C9CsX1�뮍t& � ���u�P$�����u��E    ��t��   �z������&    �H��Y��ɉX����VR��  ��농t& ���S�P$�����u��   �?����ËE���=�Et�U��.7����S��h f�f��U��WVS�u���4�E�F�]j V�r�  �EЉ4$�u$�u �u�u�u�u�uP������EЋUԃ�,�E�U��{  �u�E�V�u$�u(�u��(n �E������   �}�tD��t1�1��}�tF��8�u�E$��}�E�U��E��W�P���Eu^�E�e�[^_]� ��P;Ps��E묋C9CsX1�뮍t& � ���u�P$�����u��E    ��t��   �z������&    �H��Y��ɉX����VR�9�  ��농t& ���S�P$�����u��   �?����ËE���=�Et�U��5����S�ug f�f��U��WVS��D�] �ClP�E�P�w����{���E��E�   ��J��@t���
   �   DEȍE�u��VP���������E���  �E��P�b����MЃ���8AJ�E��l  �M��Q���}  �M�8A$��  �E��t��P�a�  �E�������E��VP�z���������  �E��E��E�    �E� �@�}��E�   t�}ȉ}Ԅ��E�F��  �}��1�   ��E��uȉE��EЍxN�@d�}����E���  1�1��}� ��  �Eԃ�0�E��}�
��  ��/�~  8]��u  �ۃ�09u���  �E�   ����  �P;P�*  ���E�����P�P;P�A  ��U�E����  1�1��}���  8���  1��E��E�P��uZ�Uą���:U���   �}(�    �}$�   �}� t�}$��}�M���]=�E��_�  �E�e�[^_]� f��Eă�P�E�P���  �E��P�E��p�p�r  ����u	�E$�    �Eą���:E΋E�v�H���f������^���������  �}��}(ҁ�   ���}$�   �G�����&    ��'    1�1��}� ��  f�1����������'    �C�<	�p����C�<��   �C�<w��ۃ�79u��^����uȋE�)�9���ރE�	ǋE���M����U�������1��}��   �u����B;B��  � �E1�8��a����U����   �]���������B;B��   � �E�������t& ��'    �ۃ�W������t& ���P�R(�E���E�������_����P;P�������    ���P�R$�����������E    �,��������������������R�P$������f����E    ������	����v ��'    �E��P�t������؋EЀx t	:X%��   �E�:X$�`������u�S�]�S�]	 �����E���)؍P���M�9u�ru�uȋU�)�9��E��	׋U��td�B;B��   ���E�����B�B;B��   � �U�E���R���1�1��}�t;8�������;����t& ��'    �U�   ��u��U�������1��}��]�uŋB;B�1  � �E1�믍�&    �Eą��  ����P�E�P��  ���E�    �7�����    ���R�P(�U���E������t��B;B�7����v ��'    ���R�P$����������E    �K�����������������8AK������E��@��   �t& ��'    8A%�z����   ��   ��    ��'    ��}(�ڀ}� E�7������t& ��'    ���R�P$����������E    �   �X����v ��'    ���R�P$�����������E    �E��c����t& ��'    �E��j P�b�  ���C����v ��'    �E��P������؋EЃ��@�M��E�    �E� �MԄ�t�M�8Y%�6  �M�8Y$�*  8YN��   �}� �  �M�8YLt	8YM��   �}�t���*  �E�    �E� �E�   �E��t�P;P��   ���P�E�����E��VP蹮������tb�E��E��E��@�F������������������}�
��:U��i����E��}���   ����   �E��{�����}��E��}��������E��P�ԭ�����}� �؋E��|   �@��������&    ���P�R(���B������������������}ԉ}������U��]-���E�e�[^_]� 1��E� �f������w����}��E��}��s����   �Q����E��@�P����E�    �E��E�   �����ËE��=�Et�U���,����S�^ f�S���\$�t$<�t$<�t$<�t$<�t$<�t$<�t$<�t$<S������4��[� f�f�f�f��S���D$�\$�L$(��R����u3���t$<�t$<Q�t$<�t$<�t$<�t$<PS������,�؃�[� �t& ���t$<�t$<Q�t$<�t$<�t$<�t$<PS�҃�,�؃�[� f�f�UWVS��,�D$X�@��   �D$�����T$���L$(Q�t$lP�t$l�t$l�t$l�t$l�t$lR�(����D$4�T$8�D$t�D$H�T$x��,����  �D$`��� �D$d�    �D$XP�D$TP�%���������  �D$\���  ��&    ��'    ����l�   P�D$(P�:����ǋ@ ���O�D$���ɉ��É�1��v ��'    �؃�8���   �D$H����  �|$L��|  �D$P���;  �D$ 1��|$T���   ��:D$�  �|$H���  �D$L����Y  ��u	�M81��8���   ��u�]83�D$�\$8��H  �ȃ�8��;  �D$H����t�P;P�  ���P�D$L�����ɺ   t;u �|$ �   ����;u�É؃�8��������1����th9w uc��t_�|$ �L$`� �=  �������t$\��B  ����'    �x;x��  �1��D$T��:D$�������͸   ���u��|$ �%  9w�  ���  �t$`�뎍t& ��'    �x;xs8��D$L�D$P���u��������G;Gsh� �D$L������    ��    �T$�L$���8P�W$������L$�T$u��D$H    �D$P���J����D$�������������������T$�L$���W�P$������L$�T$�t����D$H    ������������&    �t$`��&�t$@�D$H�T$L����V��,[^_]� �v ��'    �t$`��� tL�D$\�    ����'    �L$���P�R(���L$�������    �ɉ�t
;w u��uZ��D$`�  �D$\�    �s����v ��'    �T$�L$���8P�W$������L$�T$�����D$P    �   ������D$`�  1����������'    9w�����댋D$L�����f�f�f�f�f�f�U��WVS��D�] �ClP�E�P�w����{���E��E�   ��J��@t���
   �   DEȍE�u��VP���������E��  �E��P�b����MЃ���8AJ�E��L  �M��Q���]  �M�8A$��  �E��t��P�ay  �E�������E��VP�z��������  �E��E��E�    �E� �@�}��E�   t�}ȉ}Ԅ��E�F��  ���  ��}�f�E̋EЍxN�@d�}����E���  1�1��}� ��  �Eԃ�0�E��}�
��  ��/�g  8]��^  �ۃ�0f9u���  �E�   ����  �P;P�  ���E�����P�P;P�)  ��U�E����  1�1��}��z  8���  1��E��E�P��ub�Uą���:U���   �}(1�f��}$�   �}� t�}$��}�M���]=�E��_�3  �E�e�[^_]� �t& ��'    �Eă�P�E�P���  �E��P�E��p�p�d  ����u	�E$�    �Mą���:E�v�E�P���^�������  �E��N�����������������1�1��}� ��  f�1���������'    �C�<	������C�<��   �C�<w��ۃ�7f9u��u���f�uȸ��  )���9���ރE�	ǋE���^����U�������1��}��   ������B;B��  � �E1�8��r����U����   �]���������B;B��   � �E�������t& �ۃ�W�������t& ���P�R(�E���E�������f����P;P�������    ���P�R$�����������E    �3��������������������R�P$������m����E    ������ ����v ��'    �E��P蔣�����؋EЀx t	:X%��   �E�:X$�`������u�S�]�S�}� �����E���)؍P���M�f9u�rtf�uȺ��  )���9��E��	׋E��t]�P;P��   ���E�����P�P;P��   ��U�E���K���1�1��}�t48�������4����t& �E�   ��u��U�������1��}��]�űB;B�a  � �E1�붍�&    �Eą��F  ����P�E�P���  ���E�    �>�����    ���P�R(�E���E������t��P;P�>����v ��'    ���P�R$������"����E    �K�����������������8AK������E��@�  �t& ��'    8A%������   ��   ��    ��'    ���R�P$������*����E    �   �����v ��'    ����t*�E(�����f��E$�    �E�������&    ��'    �E��}(����1��f��E��v�����    ���R�P$�����������E    �E��:����t& ��'    �E��j P�R�  ���3����v ��'    �E��P�����؋EЃ��@�M��E�    �E� �MԄ�t�M�8Y%�6  �M�8Y$�*  8YN��   �}� �  �M�8YLt	8YM��   �}�t���*  �E�    �E� �E�   �E��t�P;P��   ���P�E�����E��VP詠������tb�E��E��E��@�6������������������}�
��:U��i����E��}���   ����   �E��{�����}��E��}��������E��P�ğ�����}� �؋E��|   �@��������&    ���P�R(���B������������������}ԉ}������U��M���E�e�[^_]� 1��E� �V������w����}��E��}��c����   �9����E��@�@����E�    �E��E�   �����ËE��=�Et�U�������S�P f�S���\$�t$<�t$<�t$<�t$<�t$<�t$<�t$<�t$<S�������4��[� f�f�f�f��S���D$�\$�L$(��R����u3���t$<�t$<Q�t$<�t$<�t$<�t$<PS������,�؃�[� �t& ���t$<�t$<Q�t$<�t$<�t$<�t$<PS�҃�,�؃�[� f�f�U��WVS��D�] �ClP�E�P�ז���{���E��E�   ��J��@t���
   �   DEȍE�u��VP�L��������E���  �E��P����MЃ���8AJ�E��<  �M��Q���M  �M�8A$��  �E��t��P��o  �E�������E��VP�ڝ��������  �E��E��E�    �E� �@�}��E�   t�}ȉ}Ԅ��E�F��  1Ҹ�����uȉE��EЍxN�@d�}����E���  1�1��}� ��  �Eԃ�0�E��}�
��  ��/�g  8]��^  �ۃ�09u���  �E�   ����  �P;P�  ���E�����P�P;P�  ��U�E����  1�1��}��s  8���  1��E��E�P��uc�Uą���:U���   �}(�    �}$�   �}� t�}$��}�M���]=�E��_�  �E�e�[^_]� �t& ��'    �Eă�P�E�P�/�  �E��P�E��p�p�
[  ����u	�E$�    �Eą���:E�v�E�H���]�������  �E��M�����������������1�1��}� �t  f�1���������'    �C�<	������C�<��   �C�<w��ۃ�79u��u����uȉ���9���ރE�	ǋE���e����U�������1��}��   ������B;B��  � �E1�8��y����U����   �]���������B;Bs}� �E��������ۃ�W�������t& ���P�R(�E���E�������n����P;P�������    ���P�R$�����������E    �;��������������������R�P$������q����E    ������0����v ��'    �E��P�������؋EЀx t	:X%��   �E�:X$�p������u�S�]�S��� �����U���)؍P���M�9u�ru�uȉ���9��E��	׋U��te�B;B��   ���E�����B�B;B��   � �U�E���S���1�1��}�t<8�������<�����    ��    �U�   ��u��U�������1��}��]�uċB;B�Q  � �E1�뮍�&    �Eą��6  ����P�E�P�5�  ���E�    �6�����    ���R�P(�U���E������t��B;B�6����v ��'    ���R�P$����������E    �K�����������������8AK������E��@�  �t& ��'    8A%������   ��   ��    ��'    ���R�P$������2����E    �   �����v ��'    ����t�E(� �����E$�    �E������E̋}(����1����E�������&    ���R�P$�����������E    �E��B����t& ��'    �E��j P���  ���S����v ��'    �E��P�d����؋EЃ��@�M��E�    �E� �MԄ�t�M�8Y%�6  �M�8Y$�*  8YN��   �}� �  �M�8YLt	8YM��   �}�t���*  �E�    �E� �E�   �E��t�P;P��   ���P�E�����E��VP�)�������tb�E��E��E��@�V������������������}�
��:U��i����E��}���   ����   �E��{�����}��E��}�������E��P�D������}� �؋E��|   �@��������&    ���P�R(���B������������������}ԉ}������U������E�e�[^_]� 1��E� �v������w����}��E��}������   �X����E��@�`����E�    �E��E�   �����ËE��=�Et�U��[����S�G f�S���\$�t$<�t$<�t$<�t$<�t$<�t$<�t$<�t$<S������4��[� f�f�f�f��S���D$�\$�L$(��R��0�u3���t$<�t$<Q�t$<�t$<�t$<�t$<PS�������,�؃�[� �t& ���t$<�t$<Q�t$<�t$<�t$<�t$<PS�҃�,�؃�[� f�f�U��WVS��D�] �ClP�E�P�W����{���E��E�   ��J��@t���
   �   DEȍE�u��VP�̔�������E���  �E��P�B����MЃ���8AJ�E��<  �M��Q���M  �M�8A$��  �E��t��P�Af  �E�������E��VP�Z���������  �E��E��E�    �E� �@�}��E�   t�}ȉ}Ԅ��E�F��  1Ҹ�����uȉE��EЍxN�@d�}����E���  1�1��}� ��  �Eԃ�0�E��}�
��  ��/�g  8]��^  �ۃ�09u���  �E�   ����  �P;P�  ���E�����P�P;P�  ��U�E����  1�1��}��s  8���  1��E��E�P��uc�Uą���:U���   �}(�    �}$�   �}� t�}$��}�M���]=�E��_�  �E�e�[^_]� �t& ��'    �Eă�P�E�P��  �E��P�E��p�p�Q  ����u	�E$�    �Eą���:E�v�E�H���]�������  �E��M�����������������1�1��}� �t  f�1���������'    �C�<	������C�<��   �C�<w��ۃ�79u��u����uȉ���9���ރE�	ǋE���e����U�������1��}��   ������B;B��  � �E1�8��y����U����   �]���������B;Bs}� �E��������ۃ�W�������t& ���P�R(�E���E�������n����P;P�������    ���P�R$�����������E    �;��������������������R�P$������q����E    ������0����v ��'    �E��P脐�����؋EЀx t	:X%��   �E�:X$�p������u�S�]�S�m� �����U���)؍P���M�9u�ru�uȉ���9��E��	׋U��te�B;B��   ���E�����B�B;B��   � �U�E���S���1�1��}�t<8�������<�����    ��    �U�   ��u��U�������1��}��]�uċB;B�Q  � �E1�뮍�&    �Eą��6  ����P�E�P��  ���E�    �6�����    ���R�P(�U���E������t��B;B�6����v ��'    ���R�P$����������E    �K�����������������8AK������E��@�  �t& ��'    8A%������   ��   ��    ��'    ���R�P$������2����E    �   �����v ��'    ����t�E(� �����E$�    �E������E̋}(����1����E�������&    ���R�P$�����������E    �E��B����t& ��'    �E��j P�R�  ���S����v ��'    �E��P�����؋EЃ��@�M��E�    �E� �MԄ�t�M�8Y%�6  �M�8Y$�*  8YN��   �}� �  �M�8YLt	8YM��   �}�t���*  �E�    �E� �E�   �E��t�P;P��   ���P�E�����E��VP詍������tb�E��E��E��@�V������������������}�
��:U��i����E��}���   ����   �E��{�����}��E��}�������E��P�Č�����}� �؋E��|   �@��������&    ���P�R(���B������������������}ԉ}������U��M���E�e�[^_]� 1��E� �v������w����}��E��}������   �X����E��@�`����E�    �E��E�   �����ËE��=�Et�U�������S�= f�S���\$�t$<�t$<�t$<�t$<�t$<�t$<�t$<�t$<S������4��[� f�f�f�f��WVS�� �\$H�t$0�D$���{���ⵃ��S�T$(R�t$\S�t$\�t$\�t$\�t$\�t$\P�����T$H�D$|�{��D$4�T$8����V��L[^_� f�f�S���D$�\$�L$(��R����u3���t$<�t$<Q�t$<�t$<�t$<�t$<PS�P�����,�؃�[� �t& ���t$<�t$<Q�t$<�t$<�t$<�t$<PS�҃�,�؃�[� f�f�U��WVS��d�] �ClP�E�P�g����ƋC���E�   ��J��@�E�t���   �
   DEЍE�}��WP�ڊ�������E��2	  �E��P�P�����8FJ���E��n  �V����  8F$�
	  �E��t��P�Y\  �E�������E��WP�r��������g  �F�E��E�    �E� �}��E�   t�}Љ}Ȅ��E�F�  �}� �E������E����t�E�    �E�   ��EЙ�E�RP�u��u��U��� �E��FN���U��E��Fd���E��+  �}� �E�    �    �E�    �.  ��&    ��'    �~ t	:^%��  :^$�  �Ë]����u�PS�2� ������  )؋MԍP���L�9M��U���  w�M�9M���  �UԋM��EЋ]��]����e�ً]��UԉE�MԋE��M��E��)��;]�r��   ;M���   �t& ��'    �M�	�E�UԃE��EЉUԋE���o  �P;P��  ���E�����P�P;P��  ��U�E���p  1�1��}��F  8��Z  1��E��E�P��us�U�����:U���   �}(�    �G    �}$�   �}� t�}$��}�M���]=�E��_��  �E�e�[^_]� �t& �E� ������&    �E���P�E�P���  �E��P�v�v�F  ����u	�E$�    �u�����:E�v�E�H���P�������  �E��@���f��}� �E�    �    �E�    �  �v 1����������'    �E�   ��������U�������1��}��]�������B;B��  � �E1�8�������E��P轆�������s����v �E�����  ����P�E�P���  ���E�    ������    ���P�R(�E���E�������b����P;P������    ���P�R$�����������E    �/������������������Eȃ�0�E��}�
��   ��/�����8]�������Ã�0�E��M�9M�r��   �M�9M���   �E�   ���  �P;P�[  ���E�����P�P;P�r  ��U�E��t1�1��}���   8��\����U����  �E���t<�Ã}�
�T����C�<	�[����C�<��   �C�<�����Ã�7�E��@�����B;B�$  � �E��밍v ��'    �UԋM��EЋ]��]����e�ً]��UԉE�MԋE��M��E��)��;]�rw;M�r�E� �M�	�E�UԃE��EЋE�Uԅ�������U���~���1��}��   �	����B;B��   � �E1��������&    �Ã�W�E��q���f����P�R(�E���E������t��P;P������v ��'    ���P�R$������|����E    �c��������������������R�P$�����������E    �����������v ��'    8FK������F�C  ��&    ��'    8F%�u����   �"  ��    ��'    ���R�P$�����������E    �   ������v ��'    ����t:�}� �E(��  � �����@����E$�    �E��F������������������u�1��}̉��}Љ�u��ك� 1ω��}���1�Eȉ�Ű}(��E�W�������t& ���R�P$�����������E    �E������t& ��'    �E��j P��  ��������v ��'    �E��P脂�����F���E�    �E� ��t	8^%����8^$�v���8^N��   �}� �c���8^Lt	8^M��   �}�t�Mȅ��  �E�    �E� �E�   �E��t�P;P��   ���P�E�����E��WP�Y�������tR�F�E��������t& �}�
��:U��y����E��}���   �Eȅ���   �E�닐�E�������&    �E��P脁�����}� ��tt�F� ����     �@   �������&    ��'    ���P�R(���B����U�����E�e�[^_]� 1��E� �(����������E��8����   ������F�����E�    �E��E�   ������ËE��=�Et�U�� ����S�e2 f�f��S���\$�t$<�t$<�t$<�t$<�t$<�t$<�t$<�t$<S�������4��[� f�f�f�f��S���D$�\$�L$(��R����u3���t$<�t$<Q�t$<�t$<�t$<�t$<PS������,�؃�[� �t& ���t$<�t$<Q�t$<�t$<�t$<�t$<PS�҃�,�؃�[� f�f�U��WVS�   ��d�] �ClP�E�P�x���E��C����J��@�E�t��f� �
   E��E�}��WP���������E���  �E��P����M�����8AJ�E��/  �M��Q���@  �M�8A$��  �E��t��P�Q  �E�������E��WP��������  �E��E��E�    �E� �@���E�   t�uĄ��E�F��  ���u��RVj�j��U��Z �E��E����U��pN�@d�u����E���  �}� �E�    �E�    �E� ��  �Eă�0�E��}�
��  ��/��  8]��w  �˃�0�u�9u�r��  �}�9}���  �E�E�����  �P;P�\  ���E�����P�P;P�s  ��U�E����  1�1��}���  8���  1��E��E�x��ul�U�����:U���   �}(�u$�    �G    �   �}� t�u$��u�M���]=�E��^��  �E�e�[^_]� ��    ��'    �E��u��PV�Ϸ  �E���V�p�p�<  ����u	�E$�    �u�����:E�v�E�H���W������Z  �E��G���f��}� �E�    �E�    �E� �,  �t& 1���������'    �C�<	�n����C��˃�W<�c����C�<w��˃�7�Q���f��}ԋE��U��uЉ����؉�����É����e��щMЉ���ڻ   9�r��   9E���   ����'    ]�ƋE׃E��uЉ}ԅ������U���M���1��}��   �4����B;B�,  � �E1�8�� ����U����   �]����r����B;Bs}� �E���]���1��y�������'    ���P�R(�E���E�������n����P;P�������    ���P�R$������{����E    �;��������������������R�P$������q����E    �����������v ��'    1�]��׃E��uЉ}ԋE���!  �P;P��  ���E�����P�P;P��  ��U�E��t1�1��}���   8�������E��P��z�����؋E��x t	:X%��   �E�:X$������}����u�SW��� ���������)��}ԉ��@���M�9}�rjw�}�9}�r`�}ԋE��U��uЉ����؉�����É����e��щMЉ���ڻ   9�����������9E������1��������&    ��'    �E�E���������U���
���1��}��]������B;B��  � �E1��������    ��'    �E����6  ����P�E�P��  ���E�    �i�����    ���P�R(�E���E�������q����P;P�i�����    ���P�R$������Q����E    �>�����������������8AK������E��@�4  �t& ��'    8A%������   �  ��    ��'    ���R�P$�����������E    �   ������v ��'    �}� t*�E(� �����@�����E$�    �E����������'    �u�1��}̉��}Љ�uȋu��ك� 1��ۉ��}(1�Eȉ�Ủ�E�W������t& ���R�P$������d����E    �E��I����t& ��'    �E��j P肭  ���,����v ��'    �E��P�x���؋E����@�M��E�    �E� �MȋM��MЄ�t�M�8Y%������M�8Y$�����8YNt�}� ������M�8YLt	8YM��   ��t�Uȅ���   �E�    �E� �   �E��t�H;H��   ���H�E�����E��WP��w������tP�E��E��@�4�����
��:M�r��E�����   �Mȅ���   �E�듍�&    �E��������&    �E��P�w�����}� ��tc�E��@�������    ��    ���P�Q(���T����U������E�e�[^_]� 1��E� �}����������E������   �����E��@�m����E�    �E��   ������ËE��=�Et�U��=�����S��' f�f�S���\$�t$<�t$<�t$<�t$<�t$<�t$<�t$<�t$<S�"�����4��[� f�f�f�f��S���D$�\$�L$(��R ��P�u3���t$<�t$<Q�t$<�t$<�t$<�t$<PS�������,�؃�[� �t& ���t$<�t$<Q�t$<�t$<�t$<�t$<PS�҃�,�؃�[� f�f���f�f�f�f�f�f�f���f�f�f�f�f�f�f���f�f�f�f�f�f�f���f�f�f�f�f�f�f���f�f�f�f�f�f�f���f�f�f�f�f�f�f�U��VS�]���C��	P��- ���{ t�C��t��P��  ���]�e�[^]�4  ����S�4  �4$�y& f�f�f�f��S���\$S�����\$ ��[�����f�f��S���\$�D$��)�RP�t$,�_� ����[�f�f�f�f�f�f�f�UW1�VS��,  ��$@  �\$ ����'    ���=   u�E ��  �@$=����   ���!  �ރ����  ���   ���   ��)���   )�����ƅ  h   RS�P� ����tƅ  ��,  [^_]ËE �@$=��u3�D$ <t؁�,  [^_]Ã�R�T$j ��$4  QSU�Ѓ� �T$둃��T$+Rj�T$5RSU���D$?�� �UW1�VS��  ��$0  �\$����'    ���=   u�E �U�@=��uS��}!�ރ���E���   ���   ��)���   )������Eh   RS�`� ����t�E��  [^_]�R��$  �T$QSU�Ѓ��T$�f�f�f�U��S����D�hDh�W��WH	��W    ��W    ��W    ��W    ��W    ��W    �|�  � X��D�$�W��W��X������WH	��W    ��W    ��W    ��W    ��W    ��W    �
�  ��W��D�$|W��W���W�����`WH	�dW    �hW    �lW    �pW    �tW    �xW    ��  �$�Y��W�`W���W�����2,  Y[h�Wh�Y�4Z    �8Z �9Z �<Z    �@Z    �DZ    �HZ    ��YL���Y`��}L  �$�Z��+  XZh�Wh�Z��Z    ��Z ��Z � [    �[    �[    �[    ��Z	��Z 	��Z    �L  �$Y�F+  Y[h`WhY�tY    �xY �yY �|Y    ��Y    ��Y    ��Y    � YL��Y`��K  �$DX��*  XZh`WhDX��X    ��X ��X ��X    ��X    ��X    ��X    �@XL��DX`�� K  ����Z�Y�Y    �tY�Y��E�]��Ã�����Y�	h�Y�-  �$��  �����DX�	hDX�i-  �$��  �����Y�	hY�H-  �$�  ������Z�	h�Z�'-  �$�  f�f�f�f�f�f�f����E�P����Et�Í�    ��    �����f�f�f�f�f����E�P�����EtÍ�    ��    U���h�Y耨���$ Y�t����$@X�h������Ã�P��  ����1�  �U��S��$�hD�E8���   ��E�J�҉�E��   ���hD��WH	h�W�4  �$�W��WH	�4  �$|W�`WH	�4  ��h    j�5�Dh W�  ��h    j�5�Dh�V�t  ��h    j�5�Dh V�Z  YXh Wh�Y�	E  XZh�Vh�Z��D  YXh VhY��D  XZh VhDX��D  �E��$�������؋]��Ð�E��X����E�� ����ÍE���P�b����$� f�f�f�f�f�U��VS�]����	S��h  �C$�$�� �H	�����]�e�[^]�t3  �������S$��R� ���H	����S�K3  �4$�3 f��S���\$S�����\$ ��[鵘��f�f��S���T$ �L$$�B��t���[Ít& �B�9�v<���B<t�r+<w��B�\$�SjQP�R�D$����[É���'    �B�)ًR�f�f�S���\$S��Z  �H	��[�f�f�f��U��WVS���]�}S�s$�Z  ���H	W�uV� �4$�� ����u�e�[^_]Í�&    ��'    �E���{,�C8S�~[  �C4�C= ���C> �C    �C    �C    �C�C�C�e�[^_]Éƃ�S�Oh  �4$�� f�f�f��U��WVS���]�}S�s$��Y  ���H	W�uV�� �4$�= ����u�e�[^_]Í�&    ��'    �E���{,�C8S��Z  �C4�C= ���C> �C    �C    �C    �C�C�C�e�[^_]Éƃ�S�g  �4$�' f�f�f���D$$�� f�f�f��D$$�� f�f�f�UWVS���\$ �D$(�l$$� �C;C��   � 1�����'    �K�s)΃�~C���E VQU�P0��C�9�q���S�P$�����uʍv ��'    ����[^_]Í�    �M;Ms(��E�C�K��9�sE���C9�s�� 농�    ���M ��PU�Q4�����uȋD$(�  ����[^_]É���'    ���S�P(������{����C�K뤍v ���1�S�P$����������T���f�f��T$�B t&�J�B��t	9�v�J��+B���������������������f�f�f�f�f��D$�@ t6�P�H��t9�w�@9�s!� Í�    ��'    �P�������'    ������f�f�f�f�f�WVS�L$�D$�Q9Qs=���t(8B�����t�A t(�r��ۉqu���Z�[^_Ð�t& ��1��Q[^_Ít& �������f�f�f�f��VS���\$ �C$�H	�P���Eu#�H	����S��.  ��$[^Ít& ��'    �H��q��ɉp�Ѓ��D$PR��  ���VS���\$ �C$�H	�P���Eu#�C���H	P�q.  �$�������$[^Ív �H��q��ɉp�Ѓ��D$PR赏  ���VS���\$ �C(�L	�C,`	�CH	�P���Eu5�C ���CH	��,P��-  ��	�$�q%  ��$[^Ít& ��'    �H��q��ɉp�����D$PR�5�  ��뫋D$�A�D$�n���f�f�f�f�f�f�f�VS���\$ �C,��	�C0�	�CH	�P���Eu5�C$���CH	��0P�_-  ��	�$��$  ��$[^Ít& ��'    �H��q��ɉp�����D$PR蕎  ��뫋D$�A�D$�n���f�f�f�f�f�f�f�VS���\$ �C(�L	�C,`	�CH	�P���Eu5�C ���CH	P��,  �C,�C,�	�$�0$  �$�8�����$[^�f��H��q��ɉp�����D$PR���  ��뫋D$�A�D$�n���f�f�f�f�f�f�f�VS���\$ �C,��	�C0�	�CH	�P���Eu5�C$���CH	P�",  �C0�C0�	�$�#  �$蘑����$[^�f��H��q��ɉp�����D$PR�U�  ��뫋D$�A�D$�n���f�f�f�f�f�f�f�VS���\$ �C0��	�C4�	�C�	�CH	�P���Eu.�C(���CH	��4P�x+  ��	�$��"  ��$[^Ít& �H��q��ɉp�Ń��D$PR赌  ��벃l$�v�����    �D$�A�D$�^���f�f�f�f�f�f�f�VS���\$ �C0��	�C4�	�C�	�CH	�P���Eu>�C(���CH	P��*  �C4�C4�	�$�9"  �$�A�����$[^Ít& ��'    �H��q��ɉp�����D$PR���  ��뢃l$�f�����    �D$�A�D$�N���f�f�f�f�f�f�f�S���\$�C�H	�C    �C    �C    �C    �C    �C    P�o�  �D$$�H	�C$F�C ��[�f�f�f�U��VS���]�U�F�B����   �J9�w:�E�j PQ�r�[�  Z�E�E�YPS�ܞ  �E���P���Eu+�e���[^]� �M�j QP�r�!�  ^�E�E�ZPS袞  �ċH��q��ɉp�ȍE��PR�Ɗ  ��붐����$RS�s�  ��룉��������E��=�Et�U��~�����=�Et�U��k~����V�� f��D$�P�H ��t";Pv-��u�P�P�PÍ�&    ��'    �Í�&    ��'    ��f�f�f�f�f�f�f�VS�T$�\$�L$�t$�D$�� �K�K�s|(~�v ��'    �����  ������ �|=���w�ȉC[^�f�f�f�f�f�f�UWVS���\$ �D$$�s$�K �n�V��σ�����9�tl$(�D$(    ���t#�t$(�C�kƅɉsu@��[^_]Ð��&    ��t��1��t$8WVRPS�)����k�k�� �k�ˍt& ��'    ��1��t$8WVRPS������� ��[^_]�f����D$�T$�P ���P$t�J�Qj RP�-�����É���'    1�Qj RP�������WVS�t$�\$�|$��t'��x#�C$j �p�C$j P�f�  ��j WVS���������[^_�U��WVS��,�]�u�C �W  ����^  �C$�K;K�@���=���?�E���8��,  ��t����C���e�[^_]Í�    �E��=�  ��   �   �}���E�FPW�7�  �C����t�S��)�RPW�=�  ���E�P�J;H��M�w�H���~���u�W���  �E���P���E�=F��   �C$��WP�M|  �C+C��P�C+CP�s$S������E���P���E�*����H��y��ɉx������E��PR�P�  ���������&    =���?��������?�����t& ��'    �e������[^_]Ív 1����������'    �M��@�    �H�� �@����ËE��=�Et�U���z����S�J f�f�f�f�f�S���D$�\$� �p�P�C$P���  ��1��C �C$t�P�Rj PS�������[�f�f��U��WVS��(�]�u�{�H	�C    �C    �C    �C    �C    �C    W�(�  �E�M���H	�C     � Q�p�P�C$P肞  ���s ���C$t$�P�Rj PS�7������e�[^_]Í�    ��    1��ۉ���ƋC$��=�Et�U��y�����H	W�B$  �4$�* f�f�f�f�f�UWVS��,�D$D�T$T�|$H�l$L�p �<$�|$@�l$���������G�����Ӊ\$�����։��É�!��|$P�É�!����Ã���!��T$�� ʈT$��   �P��u�$�\$��	���   �H��t;Hv�\$����   �H�|$P�&  �|$P�4$�|$�t$�|$�L  �|$��x8��
L$t0�H)щˉL$��9���   �$�H�|$@�t$ىH�ىw��|$��xm��
L$te�H)щ���9�}~���t$�|$ WV�p�pP�5����D$`�� �0�x�0��&    �P��u�4$�|$��	�u�|$ ������������D$@��,[^_]� ����'    �H�H������t& �9L$�v�����f��N����|$9<$�'����<������&    �p)щ���)։t$��$\$�t$�L$�L$$�\$�\$\$������    �H)щ���$\$�$�\$�L$�\$����f�f�f�f�f��UWVS���T$4�\$D�D$0�t$8�|$<�J � �����@�����̓����D$�����D$�|$ t(�J��u5��	�t/�t& ��'    ��[^_]� ��    �J��u��	�u�|$ t܋Z��t;Zv��tL�Z��xŋj)͉���9�|�9�r��|$ u:�|$ uB�T$8��T$<�P�T$@�P��[^_]� �t& �Z�Z묐��&    �J�|$ �Jt��D$��WV�r�rR������ �D$�f��U��WVS��$�u�]�F�P��N��C    �x�j �W�{�\5  ���@�V��C$�CH	�C    �C    �C    �C    �C    �C     �$��  �E�CH	�C,F���C(ZYW��H��Q��4  ���e�[^_]ÉE��W�����V��R�N�X�u���
 f�f�f�f�f�f�f�U��WVS��(�]�s0V��  ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       ��	�C0�	�C    Y_j V�=4  �C$��	�C0�	�CH	�C    �{�C    �C    �C    �C    �C     �$��  �E�CH	�C,F���C(XZWV��3  ���e�[^_]É���E��W������}�����C0�	V�P  �<$�	 f�f�f�f�U��WVS��4�u�]�F�{�P��N��C    �H�j �Q�\3  ��K$�MЉ�@�V��E�CH	�C    �C    �C    ���C    �C    �C     �Eԉ$��  �E�U���CH	�C(    � R�p�P�C,P��  ��1��E�EԉC(�C,t�P�Rj PW����XZW��P��R�2  ���e�[^_]É���E��E�ǋC,��=�Et�U��s�����CH	�u��  �����V����R�N�P�v ��W�}����Eԃ���f�f��U��WVS��8�]�s0V�{  ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       ��	�C0�	�C    Y_j V��1  �E�K$��	�C0�	�CH	�{�C    �C    ���C    �C    �C    �C     �Eԉ$�M���  �E�U���CH	�C(    � R�p�P�C,P�^�  ��1��E�EԉC(�C,t�P�Rj PW����XZWV�$1  ���e�[^_]É��/�E��B�C,��=�Et�U��q�����CH	�u��  �����C0�	V�  �<$�� ��W������}ԃ��׉�멉��f�f��WVS���t$$�\$ ���@�V��C,�CH	�P���Eu0�C$���CH	P�  �F��@�V��� [^_Ð��&    �H��y��ɉx�Ã��D$PR��|  ��밋D$���f�f�f�f�U��VS���]�U�F�B����   �J9�w:�E�j PQ�r軒  Z�E�E�YPS�<�  �E���P���Eu+�e���[^]� �M�j QP�r聒  ^�E�E�ZPS��  �ċH��q��ɉp�ȍE��PR�&|  ��붐����,RS�ӏ  ��룉��������E��=�Et�U���o�����=�Et�U���o����V�R f�VS���D$�\$� �s�p�P�C,P��  ��1��C(�C,t�P�Rj PV�������[^�U��WVS��$�u�]�F�{�H��Vىj Q��.  ���@�V��C �CH	�C    �C    �C    �C    �C    �C    �$��  �E�CH	�C(F���C$ZYW��H��Q�W.  ���e�[^_]ÉE��W�p����V��R�N�X�u��I f�f�f�f��U��WVS��(�]�s,V�[  ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       �	�C, 	Y_j V�-  �C �L	�C,`	�CH	�C    �{�C    �C    �C    �C    �C    �$���  �E�CH	�C(F���C$XZWV�H-  ���e�[^_]É���E��W�]����}�����C,�	V��  �<$�/ f�f�f�f�f�f�f��U��WVS��4�u�]�F�{�H��Vىj Q��,  ��K �MЉ�@�V��E�CH	�C    �C    �C    ���C    �C    �C    �Eԉ$��  �E�M���CH	�C$    � Q�p�P�C(P�k�  ��1��E�EԉC$�C(t�P�Rj PW����XZW��P��R�*,  ���e�[^_]É���E��E�ǋC(��=�Et�U��l�����CH	�u��  �����V����R�N�P�� ��W������Eԃ���U��WVS��8�]�s,V��
  ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       �	�C, 	Y_j V�T+  �E�K �L	�C,`	�CH	�{�C    �C    ���C    �C    �C    �C    �Eԉ$�M���  �E�U���CH	�C$    � R�p�P�C(P��  ��1��E�EԉC$�C(t�P�Rj PW����XZWV�*  ���e�[^_]É��/�E��B�C(��=�Et�U��k�����CH	�u��  �����C,�	V�  �<$�u  ��W�|����}ԃ��׉�멉��f�f�f�f�f�f�WVS���t$$�\$ ���@�V��C(�CH	�P���Eu0�C ���CH	P�  �F��@�V��� [^_Ð��&    �H��y��ɉx�Ã��D$PR�Uv  ��밋D$���f�f�f�f�U��VS���]�U�F�B����   �J9�w:�E�j PQ�r�;�  Z�E�E�YPS載  �E���P���Eu+�e���[^]� �M�j QP�r��  ^�E�E�ZPS肉  �ċH��q��ɉp�ȍE��PR�u  ��붐����(RS�S�  ��룉��������E��=�Et�U��_i�����=�Et�U��Ki����V��� f�VS���D$�\$� �s�p�P�C(P�}  ��1��C$�C(t�P�Rj PV�V�����[^�U��WVS��$�u�]�F�P��N��C    �x�j �W�?(  �F�C�@�V�D�Y_j P�#(  �F�{��@�V��F�C���@�V ��F$�CH	�C    �C    �C    �C�C(�C    �C     �C$    �$�M�  �E�CH	�C0F�C,XZW��H��Q�'  ���e�[^_]���E���V����R�N�P�� ����W����XZVS���  Y�u��r� f�U��WVS��(�]�s4V�  ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       ��	�C4�	�C    Y_j V��&  XZ�C�	�C4�	j V��&  �C(��	�C4�	�C�	�CH	�{�C    �C    �C    �C    �C     �C$    �$��  �E�CH	�C0F�C,YXWV�U&  ���e�[^_]É���E��W�j���XZhD	S���  �}�����C4�	V��  �<$�/� f�f�f�f�f�f�f��U��WVS��4�u�]�F�P��N��C    �H�j �Q��%  �F�C�@�V�D�_Zj P�%  �F�{��@�V��F�C���@�V ��F$�CH	�C    �C    �C    �C�C(�C    �C     �C$    �Eԉ$�ڽ  �E�M���CH	�C,    � Q�p�P�C0P�3�  �E����C,t6�C0�P�Rj PW�����ZYW��H��Q��$  ���e�[^_]Ít& ��'    �C01��ɉ���>�C0��=�Et�U��Ne�����CH	�u���  ����PPVS�=�  �<$�� �V����R�N�P�� �E����뢃�W�����}ԃ��f�f�U��WVS��8�]�s4V�  ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       ��	�C4�	�C    XZj V��#  _X�C�	�C4�	j V��#  �C(��	�C4�	�C�	�CH	�{�C    �C    �C    �C    �C     �C$    �Eԉ$��  �E�M���CH	�C,    � Q�p�P�C0P�h�  �E����C,�C0t(�P�Rj PW����ZYWV�2#  ���e�[^_]Í�&    1��׉�����:�C0��=�Et�U��c�����CH	�u��  ��PPhD	S�}�  �����C4�	V�z  �<$��� �E����륃�W������}ԃ��f�f�f�f�WVS���t$$�\$ ���@�V ��F$�CH	�C�C0�P���EuZ�C(���CH	P�  �F��@�V��F�C�F�C�@�V�T�F��@�V��� [^_Í�&    ��'    �H��y��ɉx�����D$PR�n  ��놋D$���f�f�f�f�U��VS���]�U�F�B ����   �J9�w:�E�j PQ�r�{�  Z�E�E�YPS���  �E���P���Eu+�e���[^]� �M�j QP�r�A�  ^�E�E�ZPS�  �ċH��q��ɉp�ȍE��PR��m  ��붐����0RS蓁  ��룉��������E��=�Et�U��a�����=�Et�U��a����V�� f�VS���D$�\$� �s�p�P�C0P��u  ��1��C,�C0t�P�Rj PV������[^�S�T$�Z$�Jd�0		�B    �B    �B    �B    ���B    �B    �B    �B     ��t& �     �@    ��9�u��Bd   �Zh��l�T$[�Ÿ  f�f����E�P����E�f�f�f�f�f�f�f�S���\$j葨  �S�@    ��T$$�P�T$(�P�C��[�f�f�f�f�f�f�f��U��WVS���}�]�E�{$�E���   �}�����   �E������p��    ��  ��u�O�P�Mz����1���    ��    �D�    ��9�u�Kd�֋Ch��~/1҉}܉u�]�v �Ћt��}�׉t���9�u�}܋u�]��t{9�tw����P謟  �����&    �E�   �E��{h�Cd�E�Ǎe�[^_]�f��C���C�Cu6�}� t�C     �e�C[^_]Ív ��'    �C    �⍴&    ��룃�h�	�_�  ��t	��P�� ��P�X�  �C�����C�Cu �}� t'�C     �C�E�诟  �E��]�����h�	�
�  �C    �׉�芟  ��S�A� �U��WVS���u�}�^��t�v ��'    ���sVW�S�����u�e�[^_]Ã�P軞  ���3�  �߃��t	��P��� ��P�w��f�f�f�f�f�VS���t$�F��t@�P�J��҉Hu3�v ���P�En������t�C�P����Su���ݍ�    ��'    �F    ��[^�f��S���\$�0		j S�����$�����Ch�S$��9�t��t��P踝  ���Ch    ��l�\$��[�.  f�f�f�f�f�f�f�S���\$S�����\$ ��[�m��f�f��S�D$�L$�\$�@�Q�%��t�Q�A+��t�#�����.�B*�Jt�J�Z��  ��t2% @  ����� ��   �Qt
��G�� [Ã�E�� [Í�    �Q�f� [�f�f��WVS�D$�|$��C�P��D$�p�9�G��t_1������'    ��t�8������9�r���7u���&    ��'    8����t��u�Q���}w8��!�[^_ø   �f�f�f����f�f�f�f�f�f�f��[l��f�f�f�f�f���D$�T$� �� ËT$�D$��f�f��U��WVS��,�E�u� �F�x����E���  �G����  �M�1����&    ���w  ������PQ�E��e� �����M�tڃ�h�   V��t  ��	��$�� ��PSV�w  ����P�Z;X�w�x���~��SV�t  ����P��=�=F�x  �E��� �@�S詙 ��PSV�v  ���   ��P�z;x�w�H���~��WV�4t  ����P��;�=F��   ��	���<W�N� ��PWV�_v  ����P�z;x�w�H���~��WV��s  ����P��=�=Fuy�E��� �@�<W��� ��PWV�
v  �������I����e��[^_]� ���������������}Ѓ�W踘 ��PWV�n  ���e��[^_]� �v ��'    �@�    �x��8 �t�����    ��'    �@�    �x��8 ������j*j�5�Ej V�k  �� �e����@�    �X�� �u�����ǍJ���Eu	��W�%� �Z��C��ۉB��PP�E�PQ�e  ����f�f�f��U��WVS��,�]�u��9���   �x���t|�J��Mԅ�tp��RP��� ����u_�O��th�E��VP�����u��$V�����}��]��1��W�;S�t\�O���E�M���   �S���Eu_�e�[^_]Í�&    �e�1�[^_]Í�    �EԋP��u���    �e��   [^_]Ív ��RSW�ߔ ������돍t& ��'    �K��y��ɉ{�����E�VR�vd  ���E��{����v ��'    �O��Q��ɉW��U����M߃��E�Q�u��=d  �]���E��4�����t!��P�� �ËE�֍P���Eu�؉��ڃ�P�_q���H��y��ɉx��PP�E�PR��c  ���Ӑ���D$��t%�?u1��w|�$��
	��t& �   �t& ��'    ��Í�    ��    �����uȃ�Ð�t& �   �ى���'    �   �ɉ���'    �   빉���'    �   멉���'    ��h<
	�3�  f����j h�
	h�E�|�  ���f�f�f�f���E��tÍ�    ��j h�
	h�E�L�  ��E���f����
	�f�f�f�f�f�U��WVS���u�N��tQ�V��t>1��
f���9^v,����t�P�z����xu���P�R����9^�Nwԅ�t��Q��  ���N��tY�F��tF1���v ��'    ��9^v,����t�P�z����xu���P�R����9^�Nwԅ�t��Q��  ���V1ۅ�tC�v ���t��P� �  �V������u��t�U�e�[^_]�ߕ  ���������������e�[^_]Ã�P���  ���w�  �N�O�����P��  ���^�  �N�������t��P�� ����P��n��f�f�f�f�f�f��S���D$���P����t
��[Ð�t& ��S�g����\$ ��[�Ze��f�f�f�f�f�WVS���\$$�D$ ��0���y����>t���[^_Í�    �D$��V�����4$�e������D$���[^_�f�f�f�f��U��WVS��(�}�]�E�W�C    ��C    �C    ��    �S��  ������G�P�n���s���C��t<1ҍ�&    �O�����C����t�A��9�u��    ��  ������F���V�dn���s��1҉C��t#��t& �O�����C����t�A��9�u��j�(n�����C1����&    ��'    �C�    ����u�1���    ��    �G�0��tF��P�!� �S���E�$�U���m���U�����C�W�u��42�40���"� ����u��e�[^_]Ã�P蟓  �$�w������on������  ��S�� f�f�f�f�f�f�f��U��WVS��,�M�]�U����  ���u��E����E��K�p��u��Q�9��"  �s��������u܉�����  ��u�G�P��l���S���ƅ�t�<�    1��K����9�u�9U�E�v���&    ��    ��9�u�E�C�M������E؉����� �C�P�l���K����t7�U�<�    �E�    �}�U�1ҍ�&    �{�<�<��;U�u�}Љ}�9M�}�v���    ��9�u�}�U܋M�s�C�҉Kt���u���  ���E؅�t��P�Α  ���E�u��@�C�4����t�P�J����Htw�E��C��t[1����&    �    ��9svB�S��    �E���t�H�y����xuϋ��P�R�}�{����빉���'    �e�[^_]Ð��&    ���P�R���x�����P�V�  ���Α  �b�����P�@�  ��踑  �}�{���[�����P�"�  �4$�ڐ  ����k����t��P�D� �����{�  ��S�2� ��P�	j��f�f�f�f��VS���L$�t$�\$���u��E����E��S����9�r �S����t�t$�D$�L$��[^������hp
	�0~  WVS�\$�|$�t$���t"�t& ��'    ����PVW�r��������u�[^_�f�f���=�E WVS�|$�\$�t$t8�G�����t��t��\$[^_�@���v ��'    �C�[^_Í�    ��h�E裕  ����t���h�E��  ���f�f�f�f�f��T$���u��E����E����f����f�f�f�f�f�f�f��D$�f�f�f�f�f���D$� �����@����� f�f�f�f�f�f��D$� �����@����� f�f�f�f�f�f�1��f�f�f�f�f�f��1��f�f�f�f�f�f��������f�f�f�f�f�������f�f�f�f�f�������f�f�f�f�f��D$� H	���D$�*���f�f�f�f�f�S���\$�C�H	P�	����\$ ��[�^��f�f�f�f�f�f�UWVS1ۃ��D$(�|$ �l$$��~!��&    �G�W)�u&��U �@4= 2uF����[^_]Í�    ��    �L$(��)�9�N��VU�P蠊 ��w9\$(~��밍�    ��RW�Ѓ����t�����9\$(��f��S���\$��@$=�1u�������[�f���S�Ѓ����t�S����S��[ÐUWVS1����D$(�\$ �l$$��~(��&    �C�S)�u&��P(�� 3uI�@$=�1uo����[^_]Ð�t& �L$(��)�9�N���WP�U��� ��{9t$(~��밍�    ��S�҃����t���9t$(�U�E ~����|�����    ��    ��S�Ѓ����t��S����S��f�f�U��WVS���]�u�{WV�g�������@=`1u(���uW�L������e��[^_]� ��    ��'    ���uS�Ѓ��ʉÃ�V������$�� f�f�f�f�f�f�f��S���D$�\$�PRS���������[� �S�D$��R��p1u[Í�    ��    [��f�f�f�f�f�f��VS���t$$�D$ �L$(�\$,��R���1u� �����@������[^� ����'    ���t$<�t$<SQVP�D$,�҃��D$��[^� f�f�f�f�f�f����L$$�D$ ��R���1u� �����@������� ��t& ���t$<�t$<�t$<�t$<QP�D$,�҃��D$��� f�f�f�f��T$��@=�1u1�Í�    ��'    ��f�f�f�f�f�f�f�S�L$�Q+Q�҉�t[Í�    ��'    ��X�Ё��1t��[��f�f�f�f�f�f�S���\$�C�S9�s���C9�vD� ��[Í�    ��    ��P(�� 3uC�@$=�1uY�������[�����������������@$=�1tۉ\$��[���v ��'    ��S�҃����t��C�S낍v ��'    ��S�Ѓ����t��C�S���C�Y����S���\$�S;Ss����S��[�f���P(�� 3u�@$=�1u�������f��\$��[�⍶    ��S�Ѓ����tًS�f�f�f�f�f�f���T$�B;Bs� Ë�H$��������1u�Í�    ��    �T$��f�f�f�f�f��D$��B ��f�f��S�T$�\$�B9Bs8X�t��H,��������1u[Í�    �H��J�@�[Ít& �ۉT$�\$[��f����T$�B9Bs�H��J�@���Ív ��H,��������1t��j�R�у��ڐS�T$�L$�B;Bs��B��[Ít& ��X4������� 2t��ɉT$�؉L$[��f�f�f�f�f�f�f��D$��B0��f�f���D$� H	�@    ���@�    �@�    �@�    �@�    �@�    �D$���  �D$�@�f�f�f�f��D$�@�f�f�f�f��D$�@�f�f�f�f��D$�T$P�f�f��D$�T$�P�T$�P�T$�P�f�f�f��D$�@�f�f�f�f��D$�@�f�f�f�f��D$�@�f�f�f�f��D$�T$P�f�f��D$�T$�P�P�T$�P�f�f�f�f�f�S���\$�C;Cs���C��[Ð�t& ��P(�� 3u#�@$=�1t߃�S�Ѓ����tуC��[�f��\$��[��f�f�f��D$�T$P�f�f��D$�T$P�f�f��T$�D$�J� H	�����H�J�H�J��H��J�H�J��H��J��H��T$�D$�;���f�f�f�f�f���D$�f�f�f�f�f���� �D$P�t$,�t$,軿����,�f�f�f���D$� �	�1����S���\$��	S�����\$ ��[�V��f�f�f�f�f�f�f���D$�    �@E��f�f�f�f�f�f�f���D$�@���f�f��D$�@�f�f�f�f����T$�D$�Jx��t�B�Bu���f������h�	�u  f�f�f�f�f�f�f��T$�D$B�D$����f�f�f�f�f�f����D$�T$	P�Pu����T`��f�f��D$�@�����f���D$�@���f�f��D$�@���f�f��D$�@���f�f���D$�@�f�f�f�f��T$�D$�P�P�T$����f�f�f�f���D$�@p�f�f�f�f��T$�L$�Bp�JpÐ�D$�@x�f�f�f�f�S���T$�D$�Zx�Bxj R���������[�f�f�f�f�f�f�f��VS���\$�{u t�Ct��[^Í�&    �s|��tD�~ t�F=�Ct�Cu��[^�f���V�w�������P�    ����tӃ�j V�҃�����m  VS���\$ �T$$�{u t�Ct�St��[^Ës|��tP�~ t�F=�Cu�St��[^�f��T$��V��������T$�H�    ����t˃�j V�у��T$��tm  f�f�WVS���D$ �T$$�L$(�X|��tk����3  ��t��[^_Ð��x �Ё���u!8�t=��3  ��[^_��������������������҉L$PRS�׃��L$�Đ�t& �����l  f�f�f��VS���D$�t$�X|��tI�{ t�����D3��[^Í�    ��S��������P������t����\$�t$��[^���~l  f�f�f�f�f�f�f�S���\$S������	�Cp    �Ct �Cu �Cx    �C|    ǃ�       ǃ�       ��[�f�f�f�VS���\$ �t$S���������tf��S�-������F|��S��������tg��S����������   ��S�<�������te��S���������   ��[^Í�    ��'    ���F|    S��������u�����'    ��ǆ�       S���������u���    ǆ�       ��[^�U��WVS�u��4�]�}�ClP�u������WSV�7�  V����XZWS������Cx����t0�X���E�SV�����YX�EԋWP�RXZWS�����4$�q������E�e�[^_]� ����Ã�V�R��������u�D����$�,� f�f�f�f�f�f�VS���\$�t$ S�M�  X�ClZPS�a���1����Ct ���Cu �Cp    �C    �sx�C��[^�f�f�f�f�U��VS�]��S�������	�Cp    �Ct �Cu �Cx    �C|    ǃ�       ǃ�       XZ�uS�]������e�[^]Éƃ�S������4$�`� UWVS��,�\$@�l$D9��  �Ed���  �s$�t$�}��t�G��j S��������Ch;D$t��t��P�  ���Ch    ��S�$����Ed���{��~0�}h1҉\$@��&    ��'    �׋\��։\���9�u�\$@�Cd�E�}u �sh�C�E�C�E�C�Ep�Cp��   �Ut�{u ��   �El���St�{lP�t$(V����XZVW�����4$�i���Y^WS����_XjS�����E�CXZ�sS��������,��[^_]Ð��&    ��    =  ������N�P�X���Ud�ƃ�1���t��t& ��    �D�    ��9�u�C$�D$������&    ��'    �s|����   �~ to�Cu�%�����    �u|����   �~ t�V=�Ut�Eu���������������������V�G�������    �@=��tȃ�j V�Ѓ���빍t& �T$��V��������T$�@=���l�����j V�Ѓ��T$�W����g  ��D$�T$��D$ �T$��   �f�f�f��D$�T$��   ËD$�T$��D$ �T$��   �f�f�f��   �f�f�f�f�f��   �f�f�f�f�f��D$+D$�T$9�G��f�f�f�f�f�f�f��   �f�f�f�f�f�U��VS�]���C�(	P�V�  �� 	���]�e�[^]�_������� 	��S�N����4$�� f�f�f�S���\$S�����\$ ��[�L��f�f��VS1����T$�\$���(	���C�.����C��[^Ã��� 	��S������4$�� f�f�f�f�f�f�S1����T$$�\$���(	���C�D$ P��  �C��[�f��D$�5
	�� �VS���\$�C����   �@.�C�5
	�5tD�@,�C�@L	�@    �@L	�@    �@L	�@     �@$L	�@(    �@,    �P0�C�P41����&    ��S�L8����u��[^Ã�jD�-�  ���@    � �	�@    �@    �@ �@ �@ �@    �@    �@    �@     �@$    �@(    �@,    �@0 �@1 �@2 �@3 �@4 �@5 �@6 �@7 �@C �C�����f�f�f�VS���\$�C����   �@.�C�5
	�5tD�@,�C�@L	�@    �@L	�@    �@L	�@     �@$L	�@(    �@,    �P0�C�P41����&    ��S�L8����u��[^Ã�jD���  ���@    � �	�@    �@    �@ �@ �@ �@    �@    �@    �@     �@$    �@(    �@,    �@0 �@1 �@2 �@3 �@4 �@5 �@6 �@7 �@C �C�����f�f�f�U��VS�]�C�( 	��t���P�R���]�e�[^]��������S������4$�� f�f�f�f�f�f�f�S���\$S�����\$ ��[�5I��f�f��U��VS�]�C�h 	��t���P�R���]�e�[^]��������S�����4$�N� f�f�f�f�f�f�f�S���\$S�����\$ ��[��H��f�f��VS���\$�t$ �C$P��  ����u��u�T$��u�C8   ����[^Ð��&    ��t�D$��~�D$�s4�C8����[^�f�WVS�\$�C,tc�{$��W�G�  ����tP�CL�s+s��tN���P�R����x8��W�J�  �ǋCL��$�R ���������[Ɖ�^_Ít& ��'    �������[^_���a  ��1��T$�J9Js���j�R�P4����������؃��f�WVS�� �\$0�t$4�C,��   �{> uR����C�{H��9C�~   �H��K�@�9���8���   ����   ����    D��� ��[^_É���'    ���j�S�P4�����t}�C4�{H����C    �C    ���C    �C> �C�C�C��L$�T$��jjj�j�SQ�P���D$#D$���t$���S�P$������T$�H����v ��'    ������� ��[^_�f�����u�{H �Ct���C=��܍�&    �C@�C�S@�CH�S�CD�C?�C�C��f�UWVS���\$ �l$$�t$(�C,���ǋCL����   ���P�R����ty����ts�{= um�{�S)��{> u�C8�H���Cс��  �   N�9�A�C��VU)�WP�C$�P�:�  �� 9�tC��)�9Ǹ    L�[^_]Í�    ��'    �t$(�l$$�\$ ��[^_]�������&    �C,u*�S4�S�S�S�C    �C    �C    �C>됍v �K8�S4���S�S�SvΉS�S�T
��S���_  f�f�f�f�UWVS��,�\$@�C,��  �{> �  �C�{H ��  �S9���  �C8�P����   CD$�CL���  ���P�R�����  �CL���P�R������  �D$�ŋKX�s\��1�)�)�9�N��{= t�C9Cu��E�;kT��  ���   �KP1ҍC$�1�1���KX�S\�D$h��  ��������������1������   C\�C\�CX�K9L$�[  ����  �l$)̓���   �����8���   �S\�   ��+CP�;CT��  ��WR�t$��  ����u��   닍C$���t$�sP�}�  ���� ����  1��C,��  �C4�C    �C    �C    �C= �C�C�C��&    ��'    �������,[^_]Ív ���(  �C,�C4�C�C�5  ŉk�C    �C    �C    �C=� ��,[^_]Í�    ��    ���j�S�P4�����t��C4�C    �C    �C    �C> �C�C�C�����v �sL�l$�6U�l$�UQ�KXQRP�C1P�sL�V�ƃ� �K���{����CP�k\�T$)�9�F��UPQ��n �CP���CX�^����1��,�������'    9C�SD�K4�CH �S���K��C@�C@�C�(�������'    ����u:����   ��h�	�b  �t& �C��������&    ������א��&    �C4���C    �C    �C    �C= �C�C�C�R�����h�	�a  ��t& ��U�K����1҅�����   �CP��t�T$�L$��P�Pq  ���T$�L$�KP�kT������v ��'    ��V�t$Q�sP�n ���KP�T$�������h�	�3a  �CL���P�R �t$���l����^�����V�t$�sXP�D$�zm ���T$�L$�X�����hL	��`  �Z  f�f�f�f�f�f�f�UWVS���D$0�t$4�l$8�xH �3  ����  �D$0�L$0�@�Q9��M  1ۋL$09�����A@�QD�y4�AH �Q�A@�y�A�D$0�P8�x,�B����   B�9��.  �D$0�@L���E  ���P�R�����  ���  �L$0�D$0�I�@�ωL$)��  �D$0�x$���    ��'    �)��&  ƃ�UVW��  �������  ��uم��  �D$0�L$0�@4�A    �A    �A    �A= �A�A�A����[^_]Ív ��'    �D$01ۀx> �������D$8� j��t$<�P4�����tI�D$0�L$0�@4�A    �A    �A    �A> �A�A�A�����t& ��UV�t$<�b�����Ã���[^_]Ív �L$0�@1ۋQ�\������)�WPV��Xk �D$@��x��������������������D$0�@,u?�D$0�L$0�@4�A�A�A�D$0�@    �@    �@    �D$0�@=����[^_]ËL$0�D$0�Q8�@4���A�A�Av��L$0�A�A�D��A�� �L$0���^��D$0�@�D$���yH �Au�޻   ������h(	�	^  �ދQ�   �g�����W  f�f���D$�xH u�P�@H�P@�P�PD�P?�P�P�P@�P��f�f��S�D$�xH t$�H1�9H�X4�HD�@H ��P@�X�H�P@�P[�f�f�f�f�f�f�f��U��WVS��(�]�s�H	�C    �C    �C    �{$�C    �C    �C    V���  ��	�C     �C ZYPW蟽  �C,    �C4    �C8    �C< �C= �C> �C? �C@    �CD    �CH �CL    �CP    �CT    �CX    �C\    �4$��������u�e�[^_]Í�&    ��'    ��V�'����CL���e�[^_]ÉE��W�-�  �H	�4$�����X�u��� f�f�f��D$$�F�  f�f�f�S���\$�{< u�C4��t��[Í�    ���s8�%F���C<�C4����f�f�f�f��S���\$�{< t�C4��t��P��k  ���C4    �C< �CP��t��P�k  ���CP    �CT    �CX    �C\    ��[�U��WVS��,�]�u�CL���  ���P�R����u`�CL���P�R �ƃ��K1�MԋKL�P����MЋ	)ԍT$�׍U�����RP�E�WP�E�P�u�u��u��Q�� ��v/����   ����$V�uS�6�  ��9����e�[^_]Í�    �U��EȍC$���EЉ։U�)�VWP��  ��9�uȋMȋŨ�t��CL�u��V�u�RWV�s�u��u�P�Q�� ��t"�u���)�VW�u�躽  ��9����e�[^_]Ã�hX	�}Z  �HT  f�f�f�f�S���\$�CL�P�R����t�C+C��[Í�    ��'    �SL�C��+C�
P�sX�sP�t$,R�Q�� CP+C\��[�f�f��UWVS��   ��$�   �D$�F9F�  �~> ��   �FL���$  ���P�Q��8D$��   �F1�D$    �|$0��$�   �D$�F$�D$��D$��~@��u;�|$ ��   �FL���L$8�QUW�t$(P�R�� ����tw��wT$,)���8�|$ t!���j�V�P4������D$�t& ��'    �D$�ļ   [^_]Ã�R�T$$W�t$$�.�  �D$$���T$9��[����t& ��'    �D$ �D$�ļ   [^_]Ít& ��'    ���j�V�P4������D$������R  UWVS���l$,�\$0�t$4�|$8�E �����E����S�u�������u����[^_]� f��C$�t$0WVP�!�  ����!у��t׋KP�E ���C= �C> �C    �C    �K\�KX�K4�C    �U�K�K�K��[^_]� �VS���\$ �t$$�C,t~�{= t<�{H ��   �C2��PS�p����L$���j jRPSQ�������D$#D$���t<�S�C�����9�s;��u���C�S���C��)�PRS�����������   ���������[^�f��S8��vH�C,��   �C4�C    �C    �C    �C�C�C���C>u'�C���C����&    ���ɈD$��   �C>����    D�����[^Ít& ��'    �C9C�SD�K4�CH ���K�S��C@�C@�C�������    �C,u*�C4�C�C�C�C    �C    �C    뉍�&    �S8�C4���C�C�CvΉC�C�D��C�\����v ��'    �C4�C�C�C�C�C�D��C����f���j�D$PS����������������UWVS��<�D$\�\$T�|$X�D$�CL��t"���P�R�D$$���� |������&    �   �D$    �D$P�k$��� �����@�����D$	��D$����U!�蕷  ���8�vT�|$`�T$�D$���D$ul��th�{> uK�{= �Q  1�1�jj j U�!�  ����!у��t���|$P��W�D$P��<[^_]� �v ��'    �CL���P�Q������   �{H t%�C9C�sD�K4�CH ���K�s��C@�C@�C�t$�L$������΍,����щ��|$ t�{= uq�D$$��j �t$lQRSP������|$l�D$@��D$D�G�D$H���G�D$P��<[^_]� ��{= uZ1�1��{> ������s+s�����������    ��    �D$�L$���D$+PS������T$�L$���������`�������D$+PS�����ǉƃ����f�f�f�VS�� �\$0�t$,�C$������F����P�͵  ����t8�{H u@�D$��j j �t$<�t$<SP�����D$ ��D$$�F�D$(���F����[^� �t& �C9C�SD�K4�CH ���K�S��C@�C@�C�f�f�f�f��WVS���t$0�\$,V�L��������!  ��V�Ȳ�����ƍS$��R��  ����u�sL��[^_Í�    �{= ��   �CL���?  ���P�R�����th�{= ��   �CL���  ���P�R������   ��t����V�P����u���T$���s,jj j SR�P�D$ #D$$������b����CL    ��[^_Ít& �{> �F����[�����{> �6�����S�=�������tċC4�C    �C    �C    �C�C�C� ���1����������'    �CL�S��+S�{P�R�S2�sXWRP�Q�S\��� 1��CX)�u�CPǉCX�{\뎍t& ����RP�sP�}^ �����K  f�f�f��S�D$�T$�H,���Ã��H4�H�HtP��~LщH��u#��t�P8��v�H4�T��H�H�P[Ð�t& �@    �@    �@    [É���'    �H�f�f�f�f�f���D$���f�f�f�f��D$,��  f�f�f��D$,���  f�f�f��D$���f�f�f�f��D$(�ֲ  f�f�f��D$(�Ʋ  f�f�f��D$���f�f�f�f��D$0馲  f�f�f��D$0閲  f�f�f�S���\$��@,    �@H P�u�����P4�@= �@> �@    �@    �@    �P�P�P��[�f�f��U��WVS��(�]�{$W�+�  ������   ���]�S���������ƋE���@,    �@H P������U�B4�B= �B> �B    �B    �B    �B�B�B�<$��  ����t����u�e��[^_]Ív ��'    �e�1�[^_]Ã�u��P�_  �<$�б  ���x:����P�_  ���`  �   �Q�����������_  �E��P�����$蜴 f�f�f�f�f�f�S���\$��	S������C$���$�α  �C�H	�\$ ��[�j���f�f�f�f�f�U��WVS��$�u�]�F�{�P��N��C    �H�j �Q��������@�V��<$�7���XZW��P��R��������e�[^_]���E��W�N����E���V����R�N�P��� �U��WVS��(�]�shV�ۼ��ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       �	�Ch 	�C    Y_j V�-����{�L	�Ch`	�<$�e���XZWV�������e�[^_]É���E��W�����}�����Ch�	V苿���<$�� f��U��WVS��$�u�]�F�{�H��Vىj Q�������@�V��<$�����XZW��H��Q�������e�[^_]���E��W������E���V����R�N�P�l� f�f�f�f�f�f�U��WVS��(�]�sdV�{���ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       ��	�Cd�	Y_j V������{��	�Cd�	�<$����XZWV�������e�[^_]É���E��W�(����}�����Cd�	V�2����<$蚱 f�f�f�f�f�U��WVS��$�u�]�F�P��N��C    �H�j �Q�?����F�C�@�V�D�_Zj P�#����F�{��@�V��F�C���@�V ��F$�C�<$�A���ZYW��H��Q��������e�[^_]��	�E�����&�V����R�N�P�԰ ��W�;����}����PPVS�9z  �<$豰 �U��WVS��(�]�slV�˹��ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       �L	�Cl`	�C    XZj V����_X�C	�Cl 	j V�����{�	�Cl4	�C 	�<$�6���ZYWV��������e�[^_]É��(�E�������W�L����}��PPh�	S�Iy  �����Cl�	V�F����<$讯 f�f�f�f�f�f�f�WVS���\$,�|$4�s$V�)�  ������   h�  W�t$,V讫  �4$��  ������   ��S�����C4����   �{,�C= �C> �C    �C�C�C�C    �C    u����[^_�f���T$��Wjj j SR�P���D$#D$���uЃ�S�B���������������������1�[^_�f�f�f���D$� �D$�����S���D$�\$��P�D$�0�CP���������t�D$    �X�\$��[�@����X�C�\$���D$��[�$���f�f�S���D$�\$��P�D$�0�CP��������t�D$    �X�\$��[������X�C�\$���D$��[�����f�f�S���\$�t$�D$�0�CP�5�������t�D$    �X�\$��[�����t& �X�C�\$���D$��[�d���f�f�S���D$�\$��P�C�t$P���������t�D$    �X�\$��[�"���f��X�C�\$���D$��[����f�f�S���D$�\$��P�C�t$P�s�������t�D$    �X�\$��[�����f��X�C�\$���D$��[����f�f�S���\$�t$�t$�CP��������t �D$    �X�\$��[�f�����    �X�C�\$���D$��[�D���f�f�U��WVS��$�u�]�F�P��N��C    �H�j �Q�����F�C�@�V�D�_Zj P�����F�{��@�V��F�C���@�V ��F$�C�<$�!���ZYW��H��Q��������u�uW�2�������t+���j �H��Q�������e�[^_]Í�&    ��'    ����P�ڋB��PR�Y������e�[^_]��	�E�����&�V����R�N�P�\� ��W������}����PPVS��t  �<$�9� f�f�f�f��U��WVS��$�u�]�F�P��N��C    �H�j �Q������F�C�@�V�D�_Zj P������F�{��@�V��F�C���@�V ��F$�C�<$�����ZYW��H��Q�����E���u�0W���������t)���j �H��Q�G������e�[^_]Í�    ��    ����P�ڋB��PR�������e�[^_]��	�E�����&�V����R�N�P�� ��W�����}����PPVS�s  �<$��� f�f�f�f��U��WVS��(�]�slV����ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       �L	�Cl`	�C    XZj V�]���_X�C	�Cl 	j V�E����{�	�Cl4	�C 	�<$�v���ZYWV�������u�uW��������t'���j �H��Q��������e�[^_]Ív ��'    ����P�ڋB��PR�������e�[^_]É��(�E�������W�8����}��PPh�	S�5r  �����Cl�	V�2����<$蚨 f�f�f�f�f�U��WVS��(�]�slV諱��ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       �L	�Cl`	�C    XZj V�����_X�C	�Cl 	j V������{�	�Cl4	�C 	�<$����ZYWV�����E���u�0W�,�������t%���j �H��Q�������e�[^_]Ð��&    ����P�ڋB��PR�Y������e�[^_]É��(�E�������W������}��PPh�	S��p  �����Cl�	V�ҳ���<$�:� f�f�f�f�f�U��WVS��$�u�]�F�{�H��Vىj Q��������@�V��<$�"���XZW��H��Q������E����P�uW�/�������t(���j �P��R�������e�[^_]Ít& ��'    ����P�ڋB��PR�Y������e�[^_]���E��W������E���V����R�N�P�S� f��U��WVS��$�u�]�F�{�H��Vىj Q�������@�V��<$�B���XZW��H��Q������E����P�E�0W�M�������t&���j �P��R�������e�[^_]É���'    ����P�ڋB��PR�y������e�[^_]���E��W� ����E���V����R�N�P�s� f��U��WVS��$�u�]�F�{�P��N��C    �H�j �Q�������@�V��<$�W���XZW��P��R������E����P�uW�d�������t���j �H��Q�������e�[^_]Ë���P�ڋB��PR�������e�[^_]���E��W� ����E���V����R�N�P蓤 f��U��WVS��$�u�]�F�{�P��N��C    �H�j �Q�<������@�V��<$�w���XZW��P��R�����E����P�E�0W��������t+���j �H��Q��������e�[^_]Í�&    ��'    ����P�ڋB��PR�������e�[^_]���E��W�0����E���V����R�N�P裣 f��U��WVS��(�]�sdV軬��ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       ��	�Cd�	Y_j V�����{��	�Cd�	�<$�L���XZWV������E����P�uW�`�������t)���j �H��Q�������e�[^_]Í�    ��    ����P�ڋB��PR�������e�[^_]É���E��W�����}�����Cd�	V�����<$耢 U��WVS��(�]�sdV蛫��ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       ��	�Cd�	Y_j V������{��	�Cd�	�<$�,���XZWV������E����P�E�0W�>�������t'���j �H��Q�������e�[^_]Ív ��'    ����P�ڋB��PR�i������e�[^_]É���E��W������}�����Cd�	V������<$�`� U��WVS��(�]�shV�{���ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       �	�Ch 	�C    Y_j V������{�L	�Ch`	�<$����XZWV�����E����P�uW��������t"���j �H��Q�p������e�[^_]Ð�t& ����P�ڋB��PR�I������e�[^_]É���E��W������}�����Ch�	V�ج���<$�@� U��WVS��(�]�shV�[���ǃ�       ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       �	�Ch 	�C    Y_j V�����{�L	�Ch`	�<$�����XZWV�����E����P�E�0W���������t ���j �H��Q�N������e�[^_]Ív ����P�ڋB��PR�)������e�[^_]É���E��W�����}�����Ch�	V踫���<$� � S���\$�CP�o�������t��[Ív ���X�C��PS��������[�f��S���\$�CP�/�������t��[Ív ���X�C��PS�{�������[�f��S���\$�CP���������t��[Ív ���X�C��PS�;�������[�f��S���\$��	S�����C$�$衛  �C�H	�$�@����\$ ��[����f��VS���t$ �\$���@�V��C�C�	P�V����C(�$�K�  �C �CH	�$�����F��@�V���[^�f�f��VS���t$ �\$���@�V��C�C�	P������C,�$��  �C$�CH	�$色���F��@�V���[^�f�f��S���\$�C��	�Cd�	�C�	P�����C(�$萚  �C �CH	��d�$�+�����	�\$ ��[阩�����&    �D$�A�D$두S���\$�C�L	�Ch`	�C�	P�+����C,�$� �  �C$�CH	��h�$軱����	�\$ ��[�(������&    �D$�A�D$두VS���t$ �\$���@�V ��F$�C�	�C�CP�����C0�$襙  �C(�CH	�$�C����F��@�V��F�C�F�C�@�V�T�F��@�V���[^�f�f�f�f�f��S���\$�C��	�Cd�	�C�	P�+����C(�$� �  �C �CH	�$辰���Cd�Cd�	�$�,����\$ ��[�/�����������������D$�A�D$끐S���\$�C�L	�Ch`	�C�	P�����C,�$蠘  �C$�CH	�$�>����Ch�Ch�	�$謧���\$ ��[������������������D$�A�D$끐S���\$�C�	�Cl4	�C 	�C�	P�$����C0�$��  �C(�CH	��l�$贯����	�\$ ��[�!�����l$뙉���'    �D$�A�D$끐S���\$�C�	�Cl4	�C 	�C�	P�����C0�$虗  �C(�CH	�$�7����Cl�Cl�	�$襦���\$ ��[������&    �l$뉉���'    �D$�A�D$�n���f�f�f�f�f�f�f��D$� �f�f�f�f���D$�T$��f�f���D$� ���f�f�f��T$�D$��� ��T$�D$�R�� f�f�f�f�f�f�f����T$�D$��R�9�w���RP�t$ hx���0  f�f�f�f����D$�����?+B�D$;D$r��Ã��t$(�/  f�f���D$�T$� �@�+D$9�G��f�f�f�f���D$�L$��   9�rR�9�����f���D$�T$�L$��t�D$�L$�T$��? ��&    ��'    ���f�f�f�f�f��D$�T$�L$��t�D$�L$�T$��? ��&    ��'    ���f�f�f�f�f��T$�L$�D$��t���T$�L$�D$�*@ �t& ��'    ��f�f�f�f�f�f���T$�D$�L$)Ѓ�t�D$�T$�L$�? ��    ��    ���f�f�f�f�f��T$�D$�L$)Ѓ�t�D$�T$�L$��> ��    ��    ���f�f�f�f�f��T$�D$�L$)Ѓ�t�D$�T$�L$�> ��    ��    ���f�f�f�f�f��T$�D$�L$)Ѓ�t�D$�T$�L$�V> ��    ��    ���f�f�f�f�f��D$+D$�f�f�f����E�f�f�f�f�f��D$� F�f�f���D$�T$��
� F�f�f�f�f�f�f���T$�D$��� ��T$�D$�R�� f�f�f�f�f�f�f��T$�D$�R�� f�f�f�f�f�f�f��T$�D$��� ��T$�D$��� ��T$�D$�R�� f�f�f�f�f�f�f��T$�D$�R�� f�f�f�f�f�f�f��T$�D$��� ��D$� �@��f�f�f��D$� �@��f�f�f�����?�f�f�f�f�f��D$� �@��f�f�f��D$� �@����Ð�D$� D$�f�f�����T$�D$��J�9�sЃ��RQPh<	�)-  f�f�f�f���D$� �f�f�f�f���D$� �P�D��f�S���L$�D$�T$�	�Y�9�wG)�9�Gڅ�tȃ�t%��SP�t$ �A< ������[Í�    ��'    � �T$�����[�SPh�	hx��,  f�f�f�f�f�f�f��S�\$�L$��B���x��x� y�@�    ��[É���'    �B�    ��f�f�f��S���\$�t$S��������[�f�f�f��S���\$�t$S��������[�f�f�f���D$� �f�f�f�f���D$� �f�f�f�f���D$� f�f�f�f��UWVS���D$0�l$<�0��V�u9T$8�����FD$8��[^_]�f�9ո����w�)�9T$8w�D$4���l$����D$8�X�D$4��ރ��D$���&    ����9�w6��8V��K���u�L$���t$�t$V�?: �����L$t���ƍ�    ������l�����    ���_���f�f�f�f�����D$� �p��t$P�t$�������f�S���\$ S�< ��P�t$S�t$�������[�f�f�f�f�f��WVS�L$������T$�D$�1�N�9�r��[^_Í�    ��'    ��)����QWR�;9 ��)��Eډ�[^_�f�f�f�f�f�f�UWVS���D$ �t$,�l$$�8������_�9�v��[^_]Í�&    )�;\$(G\$(��v �ۍC�t)�Í��VUP�9 ����u����[^_]Ð��&    �������[^_]�f�����D$� �p��t$P�t$�f������f�S���\$ S��: ��P�t$S�t$�@�����[�f�f�f�f�f��S�D$�\$�������Q��u[Í�    �B�9D$FD$�f�8�P�t��Ѓ��u�[�f�f�f�f�f�f�f��UW�����VS���t$,�\$(��t=�T$ �:�o�9�v0�t& ��'    ��V�P�t$0�7 ����u��9�w�������[^_]Ív ����[^_]�f�f�f����D$� �p��t$P�t$�v������f�S���\$ S��9 ��P�t$S�t$�P�����[�f�f�f�f�f���D$�D$����f�UWVS���D$ �|$,�l$$�0���^�t��u�������[^_]Ív ��9\$(F\$(�f��ۍC�tىÃ�W�PU��6 ����t����[^_]�f�f�f�����D$� �p��t$P�t$�v������f�S���\$ S�9 ��P�t$S�t$�P�����[�f�f�f�f�f���D$�D$����f�UWVS���D$0�t$8�l$4�|$<��C�9ƉD$r�:�v ��'    ��;t$s'��W�3PU�6 ����u����[^_]Í�&    �������[^_]�f�����D$� �p��t$P�t$�v������f�S���\$ S�68 ��P�t$S�t$�P�����[�f�f�f�f�f��WVS�T$�D$�t$��z�9�s$���8�t���    ��    8u��9�r������[^_�f�f�f�f�f��UWVS���D$ �|$$�l$,�0������^��u��[^_]Í�&    ��9\$(F\$(�f��ۍC�t)�Ã�U�PW��4 ����u����[^_]Í�&    �������[^_]�f�����D$� �p��t$P�t$�f������f�S���\$ S�7 ��P�t$S�t$�@�����[�f�f�f�f�f��S�D$�\$�������Q��u[Í�    �B�9D$FD$�f����P�t	��8t��ظ����[�f�f�f�f��VS���D$�T$� ��X�r��9�F�)�QRP�B4 ��DÃ�[^�f�f�f�f�f�f��WVS�D$�T$�L$� �X�9�w2)�9�GًL$���	�q�9��F��)�WQP��3 ����D�[^_�SRh�	hx���$  f�f��UWVS���T$0�L$4�D$8�t$@�:�_�9�wL�T$<�*�U�9�wP)�9�G�)�;T$DGT$D����9ӉT$F���PVQ�q3 �T$)Ӆ�DÃ�,[^_]�SQh�	hx��C$  RVh�	hx��2$  f�UWVS���D$,�l$0�8�_�U�Z5 ����9؉�F�)�PUW�
3 ��DÃ�[^_]�f��UWVS���T$ �t$$�D$(�*�]�9�w=)�9�G؃��t$8�5 ����9؍T5 ��F�)�P�t$4R�2 ��DÃ�[^_]�SVh�	hx��#  f�f�f�VS���D$�T$�L$�t$ � �X�9�w+)�9�Gك���9�F��)�Q�t$$P�L2 ��DÃ�[^�SRh�	hx��&#  f�f�f��T$�D$��f�f����E�f�f�f�f�f��D$�@���f�f���D$�@�����f���D$�@�����f�f��D$�@    �f�f��D$=�Eu�Ív �T$�@    ��D �f�f�f�f�f�f���D$���f�f�f�f�S���\$�D$�����?wU9ÍSv6� 9�BڍS��   v 9�s��   ���  ����?)Ӂ����?G؍S��R��<  �X�@    ��[Ã�h�	��   f�f�f�f�f�UWVS�F���\$ �l$$��t7���t$,j S�Y��������Ǎpt,�����SUV�2 �����Eu!����[^_]Í�&    ��G������'    �G    ��D �σ��t$j j �p����T$ ����f�f�f����t$ �D$ P�t$ �J����T$ �����D$�D$�2���f����f�f�f�f�f��S���H�Y��ɉX~��[Ív ��'    ��RP���������[�f�f�f�f�f�f�f�S�D$=�Eu[�f��H�Y��ɉX�[����f�f�f�f�f�f��S���D$ � �P���Eu��[Í�    �H��Y��ɉX����D$PR�E�������UWVS��,�D$@�T$L+T$H�|$D��s�C��,2)�+t$H9�w�S�����   ���\$#SPU����������t!�D$@���Q� ��   � �T$�A�
�v �@�D$��u5�D$@� �H���E�  �L$�D$@�ˉ��Fu|��,[^_]Ít& �T$@�D$H��T$L�|�����   � �륍v ��'    �D$L9D$Ht���t��D$H�|$L����u?� ��D$@���Ft���    ��    �C�    �k��+ ��,[^_]Ív ��'    ��VPS��. �D$P����C�����&    �L$��WPR�T$�w. ���L$��������VPQ�_. ���������    ��'    �p��~����x��������SQ�����������f�f�f�f�f�f��S���\$�=Ft�P���~j j j S��������@�������[�f�f�f�f�f���D$��B���x������&    ��'    ��f�f�f�f�f�f�f�VS���\$�t$��B���x��S�q�����������[^� VS���\$�t$��B���x��S�A�����������[^� VS���\$�t$��B���x��S�������R�����[^� f�f�f�f�f�f��S���\$��P���x��S��������D$��[�f�f�f�f�S���\$��P���x��S���������[�f�f�f�f�f�f�VS���t$��P�Z��P���x��V�o���������[^�f�VS���t$�\$��P�9�s�P���x��V�:���������[^�QRSh<	��  VS���\$�t$��B���x��S�������R�����[^� f�f�f�f�f�f�����D$j ��r�j P��������f�f�f�VS���\$�L$�t$��@��)�9�G�9�wj RQS���������[^�PQhF�hx��  f�f�f�f�f�WVS�|$�\$�t$+j jSW���������@��������[^_� f�f�f�f�f�f�S���T$(�L$,�D$ )�u���[� �v �D$�D$$��+j QS�t$0�'����D$4��D$���B�����ډ��[� f�f�f�f�UWVS���t$ �D$(�\$,�|$$�l$0���+J�ʁ����?9�wPSPWV���������t>��t+�����SUW�j+ ������[^_]Í�&    ��'    ������[^_]Ã�h�	��  f�f�����T$$�D$R�t$$��r�j P�R�����,�f�f�f�f�f�f�f�S���D$ �\$P�j�p�j S�#�����(��[�f�f�f�f�f�f�S���T$�D$�\$�
�I�9�w��S�t$(j PR�������([�QPh	hx��?  f�f�f�f�f�f�f��WVS�|$�t$�\$��+�D$(Pjj SW������� ��@��������[^_� f��UWVS���\$ �T$$�l$(�t$,�|$0��H��)�9�G�9�w �|$0�t$,�\$ �D$(�T$$��[^_]�2���QRh	hx��  ��T$�D$�L$�T$�T$)T$+�D$�����f�f�f�f�f����D$(�T$P�t$(j �D$,+PR�������,�f�f�f�f�f�f�WVS�\$ �|$�t$S�t$VW��������t7��t��S�t$$V�s( ����[^_ËD$� ���[^_ÐWVS�\$�t$�D$������?�J���   9�r�<
9�v��VPQj S�w����� [^_Ëz�����)�9�w1��tL��VPR��' �����F��t��B�    �r��2 �f���t���t��VPR�( ����ɐ�t& � ��뻃�h3	�
  f�f�f�f�f�S���\$�t$�t$S�*�������[�f��WVS�T$�D$�\$�t$�:�O��)�9�G�9�w��T$�t$�D$[^_�����QPh3	hx��  f�f�S���\$ S��( ��PS�t$������[�f�f�f�f�f�f�f������f�f�f�f�f��S���\$ S�( ��PS�t$�t�����[�f�f�f�f�f�f�f��UWVS���\$ �|$$�T$(�t$,��A�9��/  ����?)�9��1  9�s��VRj WS������� ��[^_]��9�w�A����Vj )�WS���e�������(Ǎ29�r$��to��VRW�.& ���؃�[^_]Í�&    9�s,��)Ճ���   ������)��u]�����y������u+� ����g�����������������������[^_]Ð��VPW�% �����3����t& ��'    ��PVW�% ���������t& ��'    ��URW�o% ���c���PWh	hx���  ��h	�  f�f�f�f�f�f�f���T$�D$+�D$�m���f�f�f�f�f�f��UWVS���T$(�D$,�l$0�\$ �t$$�:�O��)�9�G�9�w��t$$�\$ �T$,�D$(��[^_]����QPh	hx��D  f�f�S���\$$S�v& ��PS�t$�t$�������[�f�f�f�f�f�����D$� �p�P�t$�t$�������f����L$��@�P�9�wj jRQ�b������PRhF�hx��  f�f�f�f�f�f���D$=�Eu��Ð�@���f�f�f�f�WVS�\$���t$�s�D$$P���������ƍ@��t���~t-�C��RPW��# ��������Eu#[^_Í�    ��    �C���E�F���t��F    ��D [^_�f�f�f�f�f��UWVS��,�\$@�D$D�;B�t:�J��9�B���)�P�t$'VR�>�������J���Eu���,[^_]Ít& �J�����덴&    �z��o����j�ՉD$��VQ�U������D$�f�f�f�f�f�f�U����U��H�9H�w�Ít& ��'    ��j R�E������Ã�P�G&  ����&  f�f�f�f�f�f�f�UWVS���t$$�\$ ��y��t?��P�,:;h�vK��US����������P�Ѓ�t@��WQP�O" ���=Fu9����[^_]����������������x� ������&    ���ǉ���'    �@�    �h��( ��[���f�f�f�f�f��UWVS���L$$�|$(�t$ �D$,��Z�9���   )�9�G؅�tE��H�,;h�vD��UV�*����D$4�����H��ȃ�t3��SRP�! ���=Fu,����[^_]�f��x� ��̐��&    ���ԉ���'    �@�    �h��( ��SWhH	hx��  f�f�f�f�f�f�f��UWVS���\$(�t$ �|$$��tG�����?�Q�)�9���   �,;i�v=9�sY��UV�_�������Q�ʃ�u0���=FuR����[^_]Ð��&    �A���~�9�r���v ��SWR�  �����9�w���)�UV��������ϋQ��f��@�    �h��( 랃�hH	�  f���+���f�f�f�f�f��S���\$ S��! ��PS�t$������[�f�f�f�f�f�f�f�������f�f�f�f�f��S���\$ S�! ��PS�t$�������[�f�f�f�f�f�f�f��UWVS���t$$�\$ �|$(��tM�����?�B�)�9�wy�,;j�vA��US��������B�Ѓ�t8������VWP�G  ���=Fu,����[^_]�f��J�����ȍ�&    ����Սv ��'    �@�    �h��( �ă�hH	�  f��S���L$�D$�\$�=���?�R�wN9�w0r��[É���'    )�j RPQ���������[Í�    ��    ��)ЉL$�\$�D$��[�������h]	�	  f�f�f�f����j �t$�t$�n������f�f�f�f�f�WVS�\$�|$��P�r;p�w�H���~��VS���������P����=Fu[^_Í�    ��'    �@�    �p��0 [^_�f�f�f�f�f�f�f�WVS�\$�|$��B�p;r�w�J���~��VS�g�������B����=Fu��[^_Ít& ��'    �@�    �p��0 ��[^_�f�f�f�f�f�f��D$�L$�P��x=�Eu*��Í�    �D$    �L$�D$�[����t& ��'    ���P��f�f�f�f����D$$� �P��H��x���Eu5�T$ ���Ít& ��'    ��j �D$PQ� ������T$ ���Ív ���P���f�f�f�f�WVS���t$ �T$$��9�t�S��K��x@���EuX�P���Eu�����[^_�f��H��y��ɉx����D$PR��������Ӄ�j �D$PQ�p������Ë믍�&    ���S��f�f�f�f��k���f�f�f�f�f��U��WVS��8�}�]�uW�� YZ���F��U�P�RS�������u�WS�����XZVS�i������e��[^_]� �Ƌ�A�=�Et�U��D�����V�t f�f�f�f�f��U��WVS��$�]�}�u�F��@��PS�)���������VjS�����XZWS��������e��[^_]� �Ƌ�A�=�Et�U��������V�1t �U��VS���]�uS�����XZ�uS�������e���[^]� �Ƌ�A�=�Et�U��}�����V��s f�f�UWVS���t$ �D$$9�t]��)��t$,j ��P����������Ǎht-��SVU�� �����Eu7����[^_]Í�    ��'    ��G�ِ��&    ���F[��^_]Ð�G    ��D �UWVS���t$ �D$$9�tm��u��t��h�	�  ���&    ��)��t$,j ��P�=��������Ǎht ��SVU� �����Eu*����[^_]���G�損�&    ���F[��^_]Ð�G    ��D ��VS���D$$�T$(�t$,��Y��)�9�G���9�wj ʍ\$SPR�)����T$0���$[^�SRhr	hx��
  f�f�f�f�f�f�S���L$�T$�\$��@�9�w�t$RQS�{�������[� PRh�	hx���	  �VS���D$�T$�t$��Y��)�9�G���9�w�j �t$$PR�����T$ ���[^�SRhr	hx��m	  f�f�f�f�f�f��UWVS���t$ �D$$9�tm��u��t��h�	�h  ���&    ��)��t$,j ��P���������Ǎht ��SVU� �����Eu*����[^_]���G�損�&    ���F[��^_]Ð�G    ��D �ƃ��D$j �t$ �T$ �RP�F����T$ ����f�f�f�f�f�f�U��WVS��,�E�}�u� �H�9��M  ��)�;]G]��)ʁ����?9��#  9Er�9Mv(��V�uSW�u������ �e�[^_]Í�    ��    �P���ыM�ʍ89�vk�;�9M��   �E�P�E�V�uP�,����4$�u�SW�u�����U�� �J���Et��Z��s��ۉr���EԍE��PQ�~������E��o����v �U)U�VSW�u�����E�Mԃ�� �ǃ�u���E�e�[^_]É���'    ��VQW�� �E���e�[^_]Í�&    �U)2)؉E�뙃�h	�  QWh	hx��  �ËE��=�Et�U��������S�Co f�����D$(� �p�P�t$,�t$,�t$,�B�����,�f�f�f�f�f�f�f�UWVS���T$,�D$0�t$ �|$$�l$(��K��)�;T$4GT$49�w"؉l$(�|$$�t$ �T$0�D$,��[^_]�����QPh	hx��\  f�f�f�f�f�f�S���\$(S� �$S�t$,�t$,�t$,������([�f�f�f�f��D$�T$�L$)T$+�D$�s���f�����T$(�D$ �L$��r�R�T$,)�R+PQ�K�����,�f�f�f��WVS�|$�t$�\$��W�� �$W�D$,)�P+SV������ [^_�f�f�f�f�f�f���D$�T$)T$�T$�L$)T$+�D$�����f�f�f�f�f���D$�T$)T$�T$�L$)T$+�D$����f�f�f�f�f���D$�T$�L$)T$+�D$����f���D$�T$)T$�T$�L$)T$+�D$�[���f�f�f�f�f���D$�T$)T$�T$�L$)T$+�D$�+���f�f�f�f�f��S��������\$��t��S�� ���j �t$PS�$����T$ ���[�f�f�f�f�����D$j �t$ �T$ �RP������T$ ����f�f�f�f�f�f��D$�T$� 9��ËD$�T$� 9��Ã�j �t$ �t$ �t$ �
����T$ ���Ã�j �t$ �t$ �t$ �����T$ ���Ã�j �t$ �t$ �t$ �:����T$ ����S���H�Y��ɉX~��[�QQRP�q�������f�f�f�f�f�f���j��  ��� �	h0�h�	P�����f�f�f�f�f�f����j�  ��� �	h��h�	P����f�f�f�f�f�f����j�f  ��� 0	h��h	P����f�f�f�f�f�f����j�6  ���  	h0�h	P�]���f�f�f�f�f�f��U��VS�u��j��  �ÍE��P�uV�����XZVS��l  �E����=�Eu��h�h�	S� ����U�������ƃ�S�+  �4$�j �ƋE��=�Et��U�������f�f�f�f�f�U��VS�u��j�n  �ÍE��P�uV�l���XZVS�l  �E����=�Eu��h�h�	S�p����U��(�����ƃ�S�  �4$�#j �ƋE��=�Et��U��������f�f�f�f�f�U��VS�u��j��  �ÍE��P�uV�����XZVS�3l  �E����=�Eu��h0h�	S������U�������ƃ�S�  �4$�i �ƋE��=�Et��U��l�����f�f�f�f�f�U��VS�u��j�N  �ÍE��P�uV�L���XZVS��k  �E����=�Eu��hph�	S�P����U�������ƃ�S�{  �4$�i �ƋE��=�Et��U��������f�f�f�f�f�U��VS�u��j�  �ÍE��P�uV����XZVS�Sk  �E����=�Eu��h�h	S������U��x�����ƃ�S��  �4$�sh �ƋE��=�Et��U��L�����f�f�f�f�f�U��VS���]S�3 ��     �����)čE�t$PS���RV�t  �$   ��  �ÍE��PV�u�V�����XZVS�j  �E����=�Eu��h�h	S������U�������ƃ�S�)  �4$�g �ƋE��=�Et��U�������f�f�f�f�U��VS�u��j�n  �ÍE��P�uV�l���XZVS�#j  �E����=�Eu��hh$	S�p����U��(�����ƃ�S�  �4$�#g �ƋE��=�Et��U��������f�f�f�f�f�U��VS�u��j��  �ÍE��P�uV�����XZVS��i  �E����=�Eu��h`h@	S������U�������ƃ�S�  �4$�f �ƋE��=�Et��U��l�����f�f�f�f�f�U��VS�u��j�N  �ÍE��P�uV�L���XZVS�ci  �E����=�Eu��h�h`	S�P����U�������ƃ�S�{  �4$�f �ƋE��=�Et��U��������f�f�f�f�f�U��VS�u��j�  �ÍE��P�uV����XZVS��h  �E����=�Eu��h�h�	S������U��x�����ƃ�S��  �4$�se �ƋE��=�Et��U��L�����f�f�f�f�f�U��VS�u��j�.  �ÍE��P�uV�,���XZVS��)  �E����=�Eu��h��h�	S�0����U�����������S�[  �4$��d f��U��WVS��(�}j�  ���w  �Ƌ �M��WVQ�P�E�$S�jg  �E����=�Eu���p"	�{hP(h�!	S�s�����U��c����׉ƃ�S��  �4$�^d �ƋE��=�Et��U��7�����f�f��U��WVS�u��(j�  ����t  �ǍE��Ph�	V����XZVS�	f  �E����=�Eu"���E�� 	h$h� 	S�{�C�����U������ԉƃ�S�2  �4$�c �ƋE��=�Et��U������֐��j�  ��� P	h�!h8	P����f�f�f�f�f�f��U��VS��j�Q  ��XZ�uS�t   ��h �h�	S�q�������S�  �4$�.c f�f�f�f�f�f�f��D$� �	��c  �S���\$��	S��c  �\$ ��[����f�f�f�f�f�f�f��U��VS�E�u���]Ph�	V�����ZYVS�ze  �E���P���Eu�E��	�C�e�[^]Í�    �H��q��ɉp�ڍE��PR��������ȋU�ƍJ���Eu	��V�Xb �Z��C��ۉB��PP�E�PQ��������f�f�f�f�f�U��WVS��,�]����  �E���@    jP�E�P�1  ������   �}� �E��   � �u�@�tx�F;F��  � �}�E� �W��t& �����9�~K����   �~�F��)щMԉ�)�9M�NMԃ���   �ʋM9ǉF�Q��   � �����9����tW�����uO�}�   ��E��G   �늃�P�  �E�u��� p�N�F�3  �`  �E�e�[^_]Ð�t& �}� t
�u�F������uۋE�U��� P�B��PR谅���E���e�[^_]�f��M��9ǉQvP���F9�s�}� �W������t& ��'    ���V�P$�}���W��������u��=  ���e�[^_]Ë��V�P(�����uP�E�P������������V�P$���r������������P��
  �E�u��� p�N�Ft �����F�~�J������@  ��S��_ �����������&  ��S��_ f�f�f�f�f�f����	�f�f�f�f�f��D$� 0	�  �S���\$�0	S�|  �\$ ��[�/���f�f�f�f�f�f�f���D$� �	�  �S���\$��	S��  �\$ ��[�����f�f�f�f�f�f�f��UWVS���l$(;l$0�\$ t{�C�x��t����t[��    ��    ���t=������t�|$$�t,��tE � �V����
�t$<�t$<P�t$<R�Q �� ��\�������u��   ��[^_]Ít& �L$,�C�Q9�t>�8*�n�����RP�� ���   ���R���뿍t& ��'    ����E�머   �f�f�f�f�f�f��UWVS��L�l$|�Et
�D$`�@�E�D$x9D$p�D$`�X�  �D$l�@9��A  �;*t��PS�3 �����'  �D$d�T$x+T$d�D$ �D$ �D$���    ID$�D$h���D$�D$`�@�x��|$�|$`�|��C�t& ��'    ����  �D$,9���  �|$ �   ����   ���   �l$���|$���  �E��D$,    �D$0    �D$4    �D$8    �D$�D$<�������L$ht�\$p�L$� �t$D$p��t9���:\$��  ��u�|$d���  ����W��t$,�V�t$|�t$|P�t$|Q�t$|R�S�L$X�T$TU�D$,�� �˃�����։U�s  �|$ �] �������������D$,���������u~i��t�Eu^����   ����   �L$�   �   ��1Ѓ���   ����   �Ѓ����u��  ����  �u��������'    ����L$~6������g  ��   �M  ������~N����맍�    ��    ���u  ���^  �Ⱥ   ����o��������������!у���  �E     �E   �u�D$�����v ��'    ��t\�L$��������D$�������    �D$������U����ȃ��\$,�T$���D$ �] �\$0�]�������    ��'    �����Ѓ���������a�����    �D$0	E�k����t& �T$,�L$0���U �M�:  ���2  �D$`�@�D$�  �D$�-�����    �D$`�@������L$d�D$,����  D$d9D$x�z  �у��a����v ��'    �D$`�@������t$d����  \$d9\$x�V  �ɺ   �   ������D$,D$d9D$x�  ��뜋D$t�@9���   �;*�8  ��PS� ������   �D$l�@9�������t& �D$p�|$d�E �D$h���Ex4�D$pD$d9D$x�����D��E1���L[^_]Í�&    �D$�����1��|$d�u��E   �Սt& �D$�D$"D$�D$ ���������t& �D$몋D$h�E��L1�[^_]Ð��&    �T$,�M�D$�U �T$0�U��L[^_]��E     �E   �   �[�����������   ����D����ɺ   �   ����������t& ��'    �D$l;X������������&    ��'    �|$d�������T$���L$x�	��$�   ��$�   P�t$|��$�   �Q �D$,�� ���T$�	�������'    �|$d�t:�L$���D$x� ��$�   ��$�   S�t$|��$�   �P �� �ƉL$�	����ɺ   �   ������c����   �D$   �   �����UWVS��,�t$L�t$L�t$L�t$L�  �������g  �D$L�@��D$��  �D$@�t$@�@�x��t��D$���D$�   f�����t�L$H� D$H��\$�
SP�t$LR�Q������t[��t�|$u��D$��|$ �D$u��~����D$�D$L�H����   �D$L� ;D$�`  ����   �T$L�D$	B��������(  �D$�D$    �D$    �D$    �D$�F�É�����ك��L$u�L$��t��T$H������1��)�����    �L$L�D$�\$L��D$�A�L$���K�L$�K~�tt�D$@�@�_�����    ��,��[^_]Í�    �D$��t6��t1�@�I9��"����8*t�T$��QP�B� �����T$������D$L�@   뤍t& �t��D$@�@�����댍�    ��    �D$@�@�D$�����D$L�@����,[��^_]ËD$L�     �@   ��,[��^_]�f�f�f�f�f�f�f������f�f�f�f�f���F�f�f�f�f�f��F�f�f�f�f�f��D$�@��f�f�f�f�WVS�t$�������^�~Ћ�� �Լ�Ӽ����� w��v��uI�81�[^_Ð��&    �N�ɍYx&�^�h9�t�V��8�F�[^_����������������   )�����  f�S���G������t,�J0�Z4�� �Լ�Ӽ����� v�     ����0R�V ����[Ã�w�J��x��t���t!�J��[�f���u�Z���t& �J���T  f�f���������@�������f�f�f�f�f�f���f�f�f�f�f�f�f���f�f�f�f�f�f�f���	�f�f�f�f�f���	�f�f�f�f�f��{���f�f�f�f�f���k���f�f�f�f�f����f�f�f�f�f�f�f��K���f�f�f�f�f����f�f�f�f�f�f�f��+���f�f�f�f�f����f�f�f�f�f�f�f�1��f�f�f�f�f�f��1��f�f�f�f�f�f��1��f�f�f�f�f�f�������f�f�f�f�f�����D$�P�D$�H9�t+1��:*t��QR�;� ��������Í�&    ��'    �   ���f�f�f��S���D$ �\$(�$    �D$    �D$   �D$    �T�3�t$,P�R�T$1�������u
�$��   ��[�f�f�f�f��D$9D$�����D��f�f�f�f�f�f���D$� �	������S���\$��	S�����\$ ��[�����f�f�f�f�f�f�f��VS���D$�t$�P�D$�H9�t%1ۀ:*t��QR�%� ����t����[^Ð�t& �D$�F   �   �F   �����[^�f�f�f�f�f�f�f��UWVS���|$ �\$$�t$(�l$,�G�S9�t/�8*t��RP�� ����t1���v"��[^_]Ív ��'    ���   [^_]Ív ��t$(�|$$�\$ �@��[^_]��f�f�f�VS���t$ ;t$(�D$�Xt*�D$�@9�tO�;*t��PS�1� ����t9��1�[^Ð�D$$�@9�tE�;*tP��PS�� ����t/�D$�@9�u��t& �D$,�T$�0�P�@   ��1�[^Ít& �D$,�L$�H뚍v �D$;Xu���f�f����	�f�f�f�f�f��D$� �	�A����S���\$��	S�,����\$ ��[�����f�f�f�f�f�f�f��VS���T$��� ��P���������� �։��H�����t	��S��O ��S����������DP����f����T$�����f�f�����DP�����f��D$��D�f�f����D�f�f�f�f�f��D$��D�f�f����D�f�f�f�f�f����D$�8 u�x u�@�   ��Ð1���Ã�j�@   ��� x	hp�hd	P�g���f�f�f���D$�@ �f�f�f���D$�@ � �f�f�WS���D$�X`S��� ������t1��   �����B`[_Ð��   ��Gw��1ɨt�����u�������t& ��'    �   ����		�G���G�f�f�f��L$���Gr$���Os���G�������	��!�GÐ�t& ��`�L$�m� f�f�W��jP�@� ������t1��   ������_Ív ��'    �F1ɉШt�����u������v �   ��	F������@F�f���D$=@Fr5=�Gs.-@F�������Ѻ��������!F����������������D$鰲 f�f�f��S�   ���\$��D����    ��    �`  ��t�Ѓ�S�W� ����t��[Ã�j�6������ �	h��h�	P�]���f�f�f�f�f�f����	�f�f�f�f�f��D$�  	������S���\$� 	S������\$ ��[����f�f�f�f�f�f�f���D$� x	�����S���\$�x	S�����\$ ��[�?���f�f�f�f�f�f�f����jh�	j�%� ����f�f�f�f�f���jh�	j�� �j���f�f�f�f�f�UWVS��,�\$@�|$H�l$�t$L��H��@��D$    �D$    �D$    �D$    ���D$   US�t$LQWjVP�R�D$,�� ��t,�l$�����t �T$�L$!у���t����t��t1���,[^_]Ð�t& ��x�9�u�D$��,[^_]Ív ��'    ���t̋��S�t$TPVW�R ���� ��t��f�f�f�f�f�f�f���j�F������ 0	h��h	P�m���f�f�f�f�f�f����j�������  	h0�h	P�=���f�f�f�f�f�f����j�������� �"	h�)h�"	P����f�f�f�f�f�f����j�������  	h��h�	P�����f�f�f�f�f�f���D$� 	�1����S���\$�	S�����\$ ��[����f�f�f�f�f�f�f��UWVS��,�D$D�l$@�T$L�t$P�|$\�D$�D$H�]�D$�D$T�D$�D$X�D$�B9�t���*t"�T$�L$��PS�6� �����L$�T$tU;t$��   �E��|$\�|$�t$P�t$�T$L�D$@�|$X�|$�t$D�|$T�|$�|$H�A��,[^_]���v ��'    �D$�7�G�D$��xt$1�9t$���D��G��,1�[^_]Ð�|$�u��G   ��D$�@9�t&��*�a����T$��PS�o� �����T$�D����D$�G�f�f�f�UWVS���\$8�t$@�l$0�T$4�|$<9�t1�E��t$@�|$<�\$8�T$4�D$0�A ��[^_]����    ��    �E�O9�t�8*t��T$��QP��� �����T$u����   [^_]�f�f�f�f�f��UWVS���l$ �\$$�t$(�|$,WVSU�P�������t	��[^_]Ð�E��|$,�t$(�\$$�D$ �B��[^_]��f�f�f�f�f�f�f��U��VS���=�O ��   ��O�_  ���  �X1��;*�E�������ÍE�Pj j S� ���5�D��j0jh\	��� ���}� t3PP�5�DS�� ���5�DjjhJ	�� ���}� t4�0���PP�5�DV�l� �����5�Djjh,	�d� ���=� ��V�q� ��뾃�u}��P������$�R���5�D��jjhM	�� Y^�5�DS� � XZ�5�Dj
�n� ���?������ �5�Dj-jh�	��� �����������S��F ��P������� ����f�f�f�f�f�f�f����H���� ��t"�@0u� ��Í�    � ��P�����'    1���f�f�f�f�f�f���	�f�f�f�f�f��D$�  	������S���\$� 	S������\$ ��[�����f�f�f�f�f�f�f����h�U��������t��h�U����������f�f�f�f�U� U�`U��VS�E�]��C   1��C    �C`U�C U�����'    �S�K�    �    ����8u��C�U��U�U�Y��� ��Uf��U�   �    ����t�S�    ����u�jj j h S��
  ��h Sh�ES�w\��XZjh�R�)s����h�Rh�ES�V\��Y^j h�R�R   � R�	�R    �R    �R �R    �R    �R    � R    �$R �%R �dR ��R   ��R���R R�~  ��h�Rh�ES�[������R   ��R��h�Rh�ES�[������R   ��R��h�Rh�ES�][������R   ��R���QW������Rh�Rh�ES�)[�����Q   � Q�	j j h�R�Q    �Q    �Q �Q �Q �Q    �Q    �Q    � Q    �$Q    �(Q    �,Q    �0Q �1Q �2Q �3Q �4Q �5Q �6Q �7Q �CQ ��R   ��Rh 	��R Q�r����h�Rh�ES�%Z������Q   ��Q�	j j h�R��Q    ��Q    ��Q ��Q ��Q ��Q    ��Q    ��Q    ��Q    ��Q    ��Q    ��Q    ��Q ��Q ��Q ��Q ��Q ��Q ��Q ��Q ��Q ��R   ��R( 	��R�Q�p����h�Rh�ES�!Y������R   ��R�	h�Rh�ES��X������R   ��R�	h�Rh�ES��X�����P   � P���P    �P    �P    �P    �P    �P    � P    �$P    �(P    �,P    �0P    �4P    �8P    �<P    �@P    �DP    �HP    �LP    �PP    �TP    �XP    �\P    �`P    �dP    �hP    �lP    �pP    �tP    �xP    �|P    ��P    ��P    jh Ph�R��P    ��P    ��P    ��P    ��P    ��P    ��P    ��P    ��P    ��P    ��P    ��P    ��P    ��P    ��P    ��P �N'����h�Rh�ES�V������R   ��R(	h�Rh�ES�V�����|R   �xR�	hxRh�ES�mV��XZjhhR�/.����hhRh�ES�LV���s�$�E��Y���� R�s�$�E��Y���� Q�s�$�E��Y�����Q�[�$�E�Y������ P�e�[^]Ã��tq��P�> ���É�h�R�L���؉���؃��É�h�R�L���؉��뾃��É�h�R�wL���؉��뤃��É�h�R�]L���؉��늃�P�����f�f�f�f�f����jh�U������E�U��E�U���f�f�f�f����jh�U�������E�U��E�U���f�f�f�f����E��t�Ð�t& ����f�f�f�f�f��S���\$�    ��E��tI��E�;�Et*�=�U t��E� ���[�f��+��������'    � ��[Ð��&    �K����f�f�f�f������E��t$��Ph�U�fK����U��Í�    ��'    ������E��f�f�U��WVS����E�]����   �=�U t]�E�=�E�u����PV��E�K���$8	V��������u8�E�P���EuH��WS��J�����e��[^_]� ��;���뜉���'    ���u�j �rZ �E���P���Et��H��q��ɉp���E��PR蘲����뙍v �+����@����U�ƍJ���Eu	��V��; �Z��C��ۉB��PP�E�PQ�T�������f�f�f�f�f�f�f���D$�@�f�f�f�f�VS���\$ �C��	�P���Eu��S�j�����$[^Ít& �H��q��ɉp�����D$PR��������S���\$S�����\$ ��[����f�f��U��WVS���]�C��	�uP�������e�[^_]Ã��׉�S���������t	��V��: ��V�о��1��f�f�f�f�f�f��W�|$1��T$�L$�����z!�ɉB�J���J"D$�����	�B    )��B    �B    ��   ǂ      �B��1�󫍺!  ��  �B ǂ      ǂ      ���)���   ���Ƃ   _�W�|$1��T$�L$�����z!�ɉB�J���J"D$�����	�B    )��B    �B    ��   ǂ      �B��1�󫍺!  ��  �B ǂ      ǂ      ���)���   ���Ƃ   _Ã��D$ P�W ���f�f�f�f�f�f�f�VS���\$�t$9�s(�������������������R�_W �C���9�u����[^�f�f�f�f�f�f�f�����D$ P�W ���f�f�f�f�f�f�f�VS���\$�t$9�s(�������������������R��V �C���9�u����[^�f�f�f�f�f�f�f�����t$ �t$ �D� 1҅�������	�ËD$�T$�L$�T$�D$�L$�� f���D$�@�	���D$��D������'    �l$�ى���'    �D$�A�D$���S���\$�C�C�	P�D���\$ ��[黲���t& ��'    �l$�ɉ���'    �D$�A�D$뱐�D$�T$�� f��U��WVS���u�]�}�F�P��N��C    �H�W�Q�a���F�C�@�V�D�ZYWP�ra�������@�V��F�C�e�[^_]ËV����R�N�P�]7 f�f�f�f�f�f��U��WVS���]�}�sV�h@���C|    ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       �,	�C@	�C    YXWV�`��XZ�C�	�C 	WV�`����	�C�	���C�	�e�[^_]Éǃ��C�	V�&C���<$�6 f�f�f�f�f�f�f�S�T$�D$�
��I�Z��J�H�J�H�I�Z�\�J��Z�Q�[�f�f�U��VS�u�]���F�P��N��C    �H�j �Q��_���F�C�@�V�D�ZYj P��_�������@�V��F�C�e�[^]ËV����R�N�P��5 U��WVS���]�sV��>���C|    ƃ�    ƃ�    ǃ�       ǃ�       ǃ�       ǃ�       �,	�C@	�C    Y_j V�0_��XZ�C�	�C 	j V�_����	�C�	���C�	�e�[^_]Éǃ��C�	V�A���<$��4 f�f�f�f�f�f�f��VS���\$�C����   �@L	�@    �@ �@$.�C�5lD�@%,1���&    ��S�L&����$u�5pD0���t& ��S�LJ����u�C�@�	�@   �@�	�@    ��[^Ã�jh�������@    � �	�@    �@    �@ �@    �@    �@    �@     �@$ �@% �@d �C� ���f�f�f�f�f�f�U��VS�]�C����t���P�R���]�e�[^]��A������S��A���4$�3 f�f�f�f�f�f�f�S���\$S�����\$ ��[�%���f�f���D$� 	�@    ��� �	�D$��?����    ��'    �D$�A�D$���S���\$�C�	�C    �C�	P�?���\$ ��[鮭����&    ��'    �D$�A�D$뱐S�L$�D$���Y�J��L$�@    �L$B�D$[�\��f�f�f�f�f�f�f�U��WVS���]�sV��;���Cx    �C| �C} ǃ�       ǃ�       ǃ�       ǃ�       �	�C 	�C    XZ�uV�%\�����e�[^_]Éǃ��C�	V�>���<$� 2 �L$�D$���R�I��f�f�f�f�f��D$��f�f�f�f�f�S���\$��P��R�T$$����[�f�f��S���\$��P��R�T$$����[�f�f���D$�@�f�f�f�f�VS���t$��@�\|��tX�{ t$�C'P�t$�t$V�A�����[^Ít& ��'    ��S�7������P�
   ����t�j
S�҃��������f�f�f�f�f�f��S�L$�D$���Y�J��@    �D$    B�D$[��Z��f�f�f�f�f�f�f�U��WVS���]�sV��9���Cx    �C| �C} ǃ�       ǃ�       ǃ�       ǃ�       �	�C 	�C    XZj V�VZ�����e�[^_]Éǃ��C�	V��<���<$�Q0 �UWVS���D$0�|$4�\$8�D$�  ��p���V����u+�Vp��t?��R�v�������H����t2�Q����   ��1Ƀ��D$0	ʉT$4��[^_]�T���ۉ���   �Atȋqx�F;F�  �Q|� �҉$�6  �   �(����'    �F�N9���  ���F9���  � �$�J��t7����������uǋx�W�����Z����D$� ��[^_]Í�    ��1ۉD$��&    ����t����� t�=   tyw7�� ��   ��@��   �L$���t$��K �����L$��	�뵐�t& =   ti=  ��   �L$���t$�K �����L$��	��{����t& ��'    �L$���t$�7K �����L$��	��M�����    ��'    �L$���t$�K �����L$��	�������    ��'    1�	�������&    �L$���t$�K �����L$��	��������    ��'    ���V�P(�����uj�x���Q�ȹ   ���������'    ���V�P$�����t��9����v ��'    ���V�P$��Q���ыR|�T$����t��������띋F�N����������f�f��U��WVS�E߃�0�]j SP�������}� tn��E�    �P�ڋ��   ����   �zx����u��E������}ȍ}�W�}�WRj�j �u��u�PV�Q�E��,= ���})�E��M� �����f�1�E���u0�e��[^_]Í�&    =�  ~9�E��u��  ��f����E�tЋ���r��FPV�mQ�����e��[^_]ËMf��E��� �����u ��P�2������X�K�Ct3�������P��������p�ރN�Fu�y����E��L������
�ȱ���ñ���^�����S�, ���N�����S�, f�f��U��WVS�E߃�0�]j SP�������}� tW��E�    �P�ڋ��   ��tx�zx����u��E������}ȍ}�W�}�WRj�j �u��u�PV�Q�U�E��,��E���u�e��[^_]Í�&    ��'    ����J��APQ�,P�����e��[^_]��ʿ����u ��P��������X�K�Ct0�Ű����P���������p�ރN�Fu�C����o������
蕰��萰���+�����S��* ��������S��* f�U��VS�E����]�uj SP�f�������tO�}� tI�E���PV��@��tx�������t<�}� t�   ����J��APQ�=O�����e���[^]Ð��u�   �Ԑ�t& �}�����������u ��P��������X�K�Ct-软����P���������H�كI�Au�;���돉��
萯��苯���&�����S��) ��������S��) f�f�f�f�f�f��U��S�E����]�C    jSP�S������}� tZ��@�Lx�Q;Qsy����Q�C   �]��Ã�P�+�������H�كI�A��   ������&    ��'    �C��uL�   ���Z�CPS��M����������]��Ð�t& ���Q�P(������{����{�����빃���l������h�����P�������X�K�Ct	�\������
�S����N����������S�( ���������S�( U��S�E����]�C    jSP�#������}� u*�C��u�   ����J��APQ�M�����؋]��Ë�@�Lx�Q;Qs����Q�U�C   �뮐��&    ���Q�P(�����uك{�����듃�u ��P�������X�K�Ct0�l�����P��������H�كI�Au������;������
�<����7����������S�' ���������S�y' f�f�f�f��U��WVS��0�E�]�}�ƍE��C    jSP��������}� ��   �����Eԋ�@�tx�F;FrL�v ���V�P$�������;E���t@�t& �K�Q;U}1���G��F�V�C9�sa���F9�s�� �����;E���uă��������M��~� �S��uX������z��GPW�aK�����e��[^_]Ít& ���V�P(�����u/�����딐��&    1�룍�    ��    ��u��e��[^_]���F�V�Z�����u ��P��������X�K�Ct2谫����P���������p�ރN�Fu�.���1��.������
�~����y���������S��% ��������S�% f�f�f�f�f��VS���t$��@�\|��tX�{ t$�C'P�t$�t$V������[^Ít& ��'    ��S�G ������P�
   ����t�j
S�҃����轹��f�f�f�f�f�f��U��WVS�E��0�}�]�G    jWP�������}� ��   �É��Eԋ�@�\x�C;C�D  �09���   ����&    �M�Q;Q��   ��A�C�S�G9���   ���C9���   �09uԉ���u����u7�������5��P�0�������p���N�F�  �����v �G��u�   ����r��FPV� I�����e��[^_]Ív ���S�P(�����t��C�S�a����t& ���S�P$��9Eԉ������!��M�����    ��'    �M�����PQ�R4������(�������������������������S�P$������������9E��������������������P�)������x�O�Gt	�������
��������������S�6# ���o�����S�&# f�f�f�VS���t$��@�\|��tX�{ t$�C'��P�t$V�������[^Í�    ��    ��S��������P�
   ����t�j
S�҃�����-���f�f�f�f�f�f��U��S�E����]�C    jSP�3������}� u
�؋]��Ív ��@�Tx�B;Bs���B�C   �؋]��Ít& ��'    ���R�P(�����u֋���P�ڋB��PR��F����뙃�u ��P��������X�K�Ct0莧����P��������H�كI�Au�����M������
�^����Y����������S�! ���������S�! f�f�f�f�f��U��S�E���(�]�C    jSP�#������}� tz��@�Dx�P;Ps	��]��Ð���P�R$�����u����E�Z�S��RS��E���E���]��Ã�P��������X�K�CuF�<�����    ��    �����듃�uȃ�P�������X�K�Ct	�d������
�[����V����������S�  ���������S�  f�f�f�f�U��S�E����]�C    jSP�#������}� u
�؋]��Ív ����@�Dx��u�uP�R ��9E�CtӋ���P�ڋB��PR��D���؃��]��Ã�u ��P��������X�K�Ct0藥����P��������H�كI�Au�����f������
�g����b����������S� ���������S� f�f�U��S�E����]�C    jSP�3������}� tO��@�Tx�B+B��tG��~3���;EOE�R�Tx�
P�uR�Q �C���]��Ít& ��'    ���t+�C�]��Ív ���R�P������ލ�&    ��'    ����P�ڋB��PR�C���C��빃�u ��P�������X�K�Ct3�\�����P�s�������H�كI�Au������C�j������
�)����$���������S�v ��������S�f f�f�f�U��VS���]�u��C    �P�ڋB���PR�C���E���jSP��������}� tR��P�ڋBx��t1�P9Ps��:J�tB������VP�R,�����u��P�ڍt& �B����PR�B�����e���[^]Ít& ���P���u ��P�j������X�K�Ct-�3�����P�J�������H�كI�Au����뢉��
��������������S�S ��������S�C f��U��S���]��C    �P�ڋB���PR��A���E���jSP�������}� t��P�ڋBx��t5�P9Ps���P�؋]��Ë��j�P�R,�����u��P�ڍ�    �B����PR�A���؃��]��Ã�u ��P�X������X�K�Ct0�!�����P�8�������H�كI�Au�����s������
��������������S�> ���w�����S�. f�f�f�f�f�f�f�U��S�E����]jSP�������}� t1��@�Dx��t$���P�R�����t#1��]��Í�    ��    ������]��Í�    ���X�C��PS�{@����������]��Ã�u ��P�P������X�K�Ct1������P�0������X�K�Cu��������p������
���������~�����S�5 ���n�����S�% f�f��U��VS�E���]�u������C����jVP�������}� t��H���At�e���[^]� ���&    �Ax�M���jjj j PQ�R�E����E��C�E�C�e���[^]� ��u ��P�J������p�N�Ft.������P�*������p�N�Fu�����k������
����������{�����S�2 ���k�����S�" f�U��WVS��4�]��P�ڋB���PR��>���Eσ�jSP�������}� t��x���Gt�e��[^_]Ð�Gx�U���M�u�8jVQRP�EЉU܉M��u�P�W�E�#Eԃ����u�����P�ڋB��PR�T>����뤃�u ��P�1������X�K�Ct0�������P��������H�كI�Au�x����X������
�ʞ���Ş���`�����S� ���P�����S� f�f�f��U��WVS��$�]�u�}��P�ڋB���PR�=���Eۃ�jSP�{������}� t��H���At�e��[^_]Ít& ��'    �Ax�M܃��j�uWVPQ�R�E�#E������uƋ���P�ڋB��PR�4=����몃�u ��P�������X�K�Ct0�ڝ����P���������x�߃O�Gu�X����^������
誝��襝���@�����S�� ���0�����S�� f�f�f���D$� �f�f�f�f�U��WVS�]��4�E�u� p����lPS��%���$�U
���Eԉ$�,���E�u��� �@�tx�F;F��  � ��   �uԉUԋN��tQ��t& ����������u�E�e�[^_]Ð�t& �UԋB�J9��  �Uԃ��B9��N  �N� ��u���1ۉEЍ�    ��    ����t����� t�=   tiw7�� ��   ��@��   ���uЉM���3 �����M���	�븐��&    =   tI=  ub���uЉM��[3 �����M���	�념�t& ���uЉM��3 �����M���	��`������uЉM��y3 �����M���	��@���1�	��7�����&    ���uЉM��3 �����M���	������Uԃ��R�P(�����ub�E�U��� P�B��PR�:���E���e�[^_]Ív �Uԃ��R�P$�����t��K�����&    ���V�P$�����t��!����UԋB�J�f����ƃ�S�*���4$�y f�f�f�f��U��S�E����]j SP�
������}� u�؋]��Ív ��'    ��@�Lx�Q;Qs����Q�U��؋]��Ív ��'    ���Q�P(�����uً���P�ڋB��PR�9����뒃�u ��P蕿�����X�K�Ct0�^�����P�u�������H�كI�Au�ܿ���F������
�.����)����Ŀ����S�{ ��贿����S�k f�f�f�f�f�������f�f�f�f�f�������f�f�f�f�f������f�f�f�f�f������f�f�f�f�f��WVS�\$��p�ހ~u t�D$�Ft��[^_Í�&    ��'    �~|��t>� t�D$�Fu�Ft��[^_Ð��W��������@=��tՃ�j W�Ѓ����&���f�f�f��D$��J���ʋL$	J�f�f�f�f�f���D$��J�T$���!Q�f�f�f�f�f��S�T$�D$��t2��
�   t1Ƀ�������Z�ËS��	ʉS[É���'    �@   ��f�f�f�f���D$�L$��R�L�f�f�f�f�f�f�f��D$�L$��R�L�f�f�f�f�f�f�f�U��WVS�E��0�]j SP�h������}� tM��E�    �x�ߋ��   ����tf�
���wx�u������M̍M�Q�M�P�E�j�j WVRP�Q��,�E��u�e��[^_]Ð��&    ����z��GPW�7�����e��[^_]�誦����u ��P�ܼ�����X�K�Ct0襗����P輼������x�߃O�Gu�#����u������
�u����p���������S�� ���������S� f������f�f�f�f�f��U��WVS�E��0�]j SP�8������}� tM��E�    �x�ߋ��   ����tf�
���wx�u������M̍M�Q�M�P�E�j�j WVRP�Q��,�E��u�e��[^_]Ð��&    ����z��GPW��5�����e��[^_]��z�����u ��P謻�����X�K�Ct0�u�����P茻������x�߃O�Gu�����u������
�E����@����ۻ����S� ���˻����S� f������f�f�f�f�f��U��WVS�E��0�]j SP�������}� tM��E�    �x�ߋ��   ����tf�
���wx�u������M̍M�Q�M�P�E�j�j WVRP�Q��,�E��u�e��[^_]Ð��&    ����z��GPW�4�����e��[^_]��J�����u ��P�|������X�K�Ct0�E�����P�\�������x�߃O�Gu�ú���u������
��������諺����S�b ��蛺����S�R f������f�f�f�f�f��U��WVS�E��0�]j SP��������}� tM��E�    �x�ߋ��   ����tf�
���wx�u������M̍M�Q�M�P�E�j�j WVRP�Q��,�E��u�e��[^_]Ð��&    ����z��GPW�|3�����e��[^_]�������u ��P�L������X�K�Ct0������P�,�������x�߃O�Gu蓹���u������
����������{�����S�2 ���k�����S�" f������f�f�f�f�f��U��WVS�E��0�]j SP�������}� tM��E�    �x�ߋ��   ����tf�
���wx�u������M̍M�Q�M�P�E�j�j WVRP�Q��,�E��u�e��[^_]Ð��&    ����z��GPW�L2�����e��[^_]�������u ��P�������X�K�Ct0������P���������x�߃O�Gu�c����u������
赒��谒���K�����S� ���;�����S�� f������f�f�f�f�f��U��WVS�E��0�]j SP�x������}� tM��E�    �x�ߋ��   ����tf�
���wx�u������M̍M�Q�M�P�E�j�j WVRP�Q��,�E��u�e��[^_]Ð��&    ����z��GPW�1�����e��[^_]�躠����u ��P�������X�K�Ct0赑����P�̶������x�߃O�Gu�3����u������
腑��耑��������S�� ��������S�� f������f�f�f�f�f��U��WVS�E��0�]j SP�H������}� tM��E�    �x�ߋ��   ����tf�
���wx�u������M̍M�Q�M�P�E�j�j WVRP�Q ��,�E��u�e��[^_]Ð��&    ����z��GPW��/�����e��[^_]�芟����u ��P輵�����X�K�Ct0腐����P蜵������x�߃O�Gu�����u������
�U����P���������S�
 ���۵����S�
 f������f�f�f�f�f��U��WVS�E��0�]j SP�������}� tM��E�    �x�ߋ��   ����tf�
���wx�u������M̍M�Q�M�P�E�j�j WVRP�Q$��,�E��u�e��[^_]Ð��&    ����z��GPW�.�����e��[^_]��Z�����u ��P茴�����X�K�Ct0�U�����P�l�������x�߃O�Gu�Ӵ���u������
�%���� ���軴����S�r	 ��諴����S�b	 f������f�f�f�f�f��U��WVS�E��0�]j SP��������}� tM��E�    �x�ߋ��   ����tf�
���wx�u������M̍M�Q�M�P�E�j�j WVRP�Q(��,�E��u�e��[^_]Ð��&    ����z��GPW�-�����e��[^_]��*�����u ��P�\������X�K�Ct0�%�����P�<�������x�߃O�Gu裳���u������
����������苳����S�B ���{�����S�2 f������f�f�f�f�f��U��WVS�E��0�]j SP�������}� tM��E�    �x�ߋ��   ����tf�
���wx�u������M̍M�Q�M�P�E�j�j WVRP�Q,��,�E��u�e��[^_]Ð��&    ����z��GPW�\,�����e��[^_]��������u ��P�,������X�K�Ct0�������P��������x�߃O�Gu�s����u������
�Ō��������[�����S� ���K�����S� f������f�f�f�f�f��U��WVS�E��0�]j SP�������}� tM��E�    �x�ߋ��   ����tf�
���wx�u������M̍M�Q�M�P�E�j�j WVRP�Q0��,�E��u�e��[^_]Ð��&    ����z��GPW�,+�����e��[^_]��ʚ����u ��P��������X�K�Ct0�ŋ����P�ܰ������x�߃O�Gu�C����u������
蕋��萋���+�����S�� ��������S�� f������f�f�f�f�f��VS�� �\$,�t$�C   �C    ��l�C�  V����XZVS�����4$�����$[^�f�f�f�f�f�f�f�WVS�t$�\$���~lWS���XZ�t$ W���Y_jV�������[^_� f�f�f��UW��VS�Ɖ�e�-    ���L$���    )�t!Ã�WSV襰 �����u������| t�D$��[^)�_]�f�f�f�f�f�f���D$�     �@ ÐWVS�|$�\$��tQ���uKe�5    �����1��    ��t& ������<u%���R�i� ����u�;�C ��[^_Í�&    [1�^_�f�f�f�f�f�U��S���E�]��=����;w���	��t���t1ۉ؋]��Í�&    ��'    ��P�u�� �����tԋU�C��u�j jj P薟 �؃��]��Ã�t	��P�� ��P裇��f��S���T$�\$��=����;w���	��t���t��1�[Ð��P�t$ �֓ �����t��C����[�f�f�f�f�f�f�f���D$� �����f�f�U����E�0艓 ���Ã�t	��P�- ��P����f�f��D$� �f�f�f�f��VS���\$���tW�{ t8e�5    ������    ���    ������<u%���R誎 ����u��    ����[^Ð�t& �    ��1�[^�f�����f�f�f�f�f��UWVSe�-    ���|$ �t$$�\$(��t& �������| u��W�
�����SVP�� �����t׃�[^_]�f�f�f�f�f�f�f��VS���\$ �t$$�t$����������[^�����f�f�f�f�f�f�VS1ۃ��t$��u1���t$�������L$ �T$������É�[^Ít& ��'    ���t$�d������T$���v���9Ɖ�t�����[^�f�f�f�f�U��WV�}�u���u�*������uWVP腫 ���e�^_]Ã�t	��P�T ��P�+���f�f�f�f�f���D$� �D$� � �VS��P�t$\V�����ZY�T$RP�Y� ��1҅�u#�\$$��V������jj j P�� )Ã��ڃ�D��[^�S���\$�t$,S變������[� f�f���D$�@�f�f�f�f��D$�@�f�f�f�f�VS���\$ �C��	�P���Eu��S�Z�����$[^Ít& �H��q��ɉp�����D$PR��v�����͋D$� �	�����S���\$��	S�����\$ ��[�z��f�f�f�f�f�f�f���D$� �	�a����S���\$��	S�L����\$ ��[�z��f�f�f�f�f�f�f���D$� �	�!����S���\$��	S�����\$ ��[�?z��f�f�f�f�f�f�f���D$� �	������S���\$��	S������\$ ��[��y��f�f�f�f�f�f�f��S���\$S�����\$ ��[��y��f�f��VS���\$ �C�	�P���Eu��S������$[^Ít& �H��q��ɉp�����D$PR�eu�����͋D$� (	�����S���\$�(	S�����\$ ��[�Oy��f�f�f�f�f�f�f���D$� @	�a����S���\$�@	S�L����\$ ��[�y��f�f�f�f�f�f�f���D$� X	�!����S���\$�X	S�����\$ ��[��x��f�f�f�f�f�f�f��S���\$S������\$ ��[�x��f�f��U��VS�]���C��	�uP�Ç�����e�[^]Ã���S让���4$���  f�f�f�S���\$�t$S������	��[�f��S���\$�t$S������	��[�f��S���\$�t$S�n�����	��[�f��S���\$�t$S�N�����	��[�f��U��VS�]���C�	�uP�������e�[^]Ã���S�����4$��  f�f�f�S���\$�t$S�����(	��[�f��S���\$�t$S�����@	��[�f��S���\$�t$S�n����X	��[�f��U��WVS��$j j � �$���x� �X�$�)�������SWP薣 XZhz	j � Y�E�[P�u蚢 �E����E�;Et�8 t[���	��&    �؋E�     �E�    ��v ��'    �؍�&    ��'    ��Vj �$ �4$�m������e�[^_]�f���	������w
��	��v����ɡ�	�M����G�	��E�    뤃�t	��P��  ��P�m��f�f�f�f�f�f��U��WVS��$j j � �$���X� �X�$�	�������SWP�v� XZhz	j �m Y�E�[P�u�G� �E����E�;Et�8 t[���	��&    �؋E����E�    ���    ��    �؍�&    ��'    ��Vj � �4$�M������e�[^_]�f�� 	������w
�	��v���������v�E� 	��E�    먐��&    �E�	�����t	��P�e�  ��P�<~��f�f�f�f�f�f�U��WVS��$�M�Ej j �u�M܉E��^ �$���� �X�$��~�����E�SWP�6� XZhz	j �- ��Vhd	�u���� ������v2�.�- 	������vb��������vl�- 	�>�E��    �%��t& �E����>�    ���؍�&    ��'    �]��Sj � �]���e�[^_]�����-	��v���������w��-	�>뒃�t	��P�D�  ��P�}��f�f�f�f�f��WV�z	�   ���D$�t$�     �u��^_Ã�h�	�l���f�f�f�f�f�f��D$�     �f�f��1��f�f�f�f�f�f��1��f�f�f�f�f�f��U��WVS��$�}j j �� �$��蕡 �X�$�F}�����E�SVP貟 �E[^�pj � ���u�u�uW�ϡ ��XZ�u�j � Y�u��Т������u� �e�[^_]Ã�t	��P�0�  ��P�|��f�f�f��S���\$�C����  �@`��@`��@o��@o��@L	�@L	�@ 0	�@$3	�@(L	�@,6	�@0=	�@4D	�@8L	�@<V	�@@_	�@Df	�@Ho	�@Ls	�@Pw	�@T{	�@X	�@\�	�@`�	�@d�	�@h�	�@l�	�@p�	�@t�	�@x�	�@|�	ǀ�   �	ǀ�   �	ǀ�   �	ǀ�   �	ǀ�   �	ǀ�   �	ǀ�   �	ǀ�   �	ǀ�   �	ǀ�   �	ǀ�   �	ǀ�   �	ǀ�   �	ǀ�   �	ǀ�   	ǀ�   	ǀ�   		��[Í�    ��    ��h�   �������@    � ���@    �@    �@    �@    �@    �@    �@     �@$    �@(    �@,    �@0    �@4    �@8    �@<    �@@    �@D    �@H    �@L    �@P    �@T    �@X    �@\    �@`    �@d    �@h    �@l    �@p    �@t    �@x    �@|    ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ǀ�       ƀ�    �C�����f�f�f�f��	�f�f�f�f�f��D$� P	鑠���S���\$�P	S�|����\$ ��[�/o��f�f�f�f�f�f�f��U�   ��WVS��|����\	��   �U�E󥍵|���)Ѝ��   �X�����t���)̹   �\$���������f��N�O�KkPRQ�?� ��t����Dj �$����f�U1҉�VS�E��0�\$��jj����5lDRP�CP�$0���� ;E��w*)Ã��CVP�u�� ���e���[^]Í�    ��    �������f�f�f�f��UWVS���L$ �D$$�t$(�|������t& ��������tq9���   <%��u��N��st��ztu1���%����ɉ���'    �D$,����u��9���   �����C����u����D$,��u�����'    � ��+D$ ��[^_]����������������~u���T����D$,���h�D$0�0��)�PS��������~Ã��l$,�,����t& ��S�t$,����f����	�f�f�f�f�f��D$� � 	�  �S���\$�� 	S��  �\$ ��[��l��f�f�f�f�f�f�f���D$� � 	�����S���\$�� 	S�l����\$ ��[�l��f�f�f�f�f�f�f��U��WVS��,�E�H�@��R���%��   ���E�F��   ~+����   ����   �E��jh�	P�fp����t& ��u{�E��jh�	P�Hp���E���P���EtG�H��Y��ɉX�:�M���E�QR��g�����E��"f��]��PQS�ҋE���P���Eu��t& �e�[^_]Ð��&    �E��jh% 	P��o��냍t& ��'    �E��jh 	P�o���`������&    �E��jh�	P�o���@����U�ǍJ���Eu	��W��  �Z��s��ۉr��U�PPRQ�g�����ِU��WVS���E�]���F��   ~P��t+��uv��jh�	S�o�����e��[^_]� ��&    ��jh 	S��n�����e��[^_]� ���u+��jh�	S��n�����e��[^_]� ��    ��    ��jh% 	S�n�����e��[^_]� ���jh�	S�n�����e��[^_]� ��ǍJ���Eu	��W��  �Z��s��ۉr��U�PPRQ��e������f�f�f�f�f���=[ t��DÐ��h[�ß������t'��h[������h`Dh�Dh�#�B ����D���f�f�f�f�f�f��� 	�f�f�f�f�f��� 	�f�f�f�f�f��D$�T$��T$�P� f�f�f�f�f�f��T$1��L$9Jt�����������������D$9���f�f�f���f�f�f�f�f�f�f���f�f�f�f�f�f�f��i��f�f�f�f�f����h��f�f�f�f�f��S��$�\$,�t$4�)� ���T$RPS�0�����(��[� f�f�f��S��$�\$,�t$4��� ���T$RPS� �����(��[� f�f�f���D$� p"	�����S���\$�p"	S�����\$ ��[�_h��f�f�f�f�f�f�f��VS���D$ �\$(�t$$��J��`'u1�9St'��[^Ív �D$��VRP��1��T$�t$��9Su�;3����[^�f�f�f����f�f�f�f�f�f�f���g��f�f�f�f�f����D�f�f�f�f�f���D�f�f�f�f�f�S���L$$�D$ �Q�	��[��`'u��P��[� ��    ��QRP�D$�Ӄ��D$��[� f�f�f��D$�[�f�f���[�f�f�f�f�f��}"	�f�f�f�f�f��D$� �"	�����S���\$��"	S������\$ ��[��f��f�f�f�f�f�f�f����Kw{UWV��S�$� #	��&    ��'    ��tL�^1�;^}"�n�<[���^�|� ��t�D$��O�G��[^_]Ít& ��'    ��t�D$��u��t& 1��܍�    ��    1�Í�    ��'    WVS�X;X}5�p�<[���X�4����Å����u��t�    �V���N[^_�f�[1�^_Ív ��'    UW��VS�Ë@�ω�� �F��    ��    ��uB<K��   �C��҃C0�����j 1ɉ���������ZtO�p�C� <r��<V��u��C��t��҃C0	����������t���҃C0	�����몍t& ��'    [1�^_]É���'    ��uL<FuH9�u�Bf���tK��u�E    ��9�t(�m �E ��u��E    ��9�u���������������[��^_]É���'    �E    븍�&    VS�Ës�����R����Ot	��u5[^�f���u,�C0�    j �����s�������Z[^Í�&    ��'    �C0�   �Ґ�t& �H�9St1�Ð�t& UWVS�Y���X�y uM1ۋH��������8�s�P���C�����ɺ -	f�:��   �����-	u�1���[^_]Ív �Y�X�Y�KЀ�	v	��_�/  ��_�|   �K�1Ҁ�	w-f��ҍL��9�w��P�: t-�Z�X���_t/�ʍKЀ�	vՍK���w��ҍL���ˍt& 1ۉ��ݍv ��'    ��;H �g����@(�@����[^_]�f�1��ߋr���t$��   �X�h�z�$    9�|$}*�p�<[���X�<���t�t$�   �<$�w�t$�w�4$�p,��tC�J�rp09�������P�<[���X����������   �J�Љr�����h�X빋J�r뻍K���������Z�����t& ��W��V��S��t�v �;Kw��$�0$	f��[��u�[^_Ð�t& �[��t& ��'    �K�9u��K���������[�Ǎt& ��K�損�&    S����   ���   t�Y��   ���  ��[Í�&    �T$��ƀ�    ��  h�   �   P�D$��  �D$��1ɋT$��   릐UW1�V��S� 1����ntL�B�1�<	w*�1ۍH��    ��    ������\B��Q��B�<	v�1�;[^_]����������������Pf� �������P렍�    ��    �P;P}HS�H�R���P����t$�@   ���V����C��[���������������1�[Í�    ��    1�Í�    ��'    S�P���<_t#<nt�C�����S�:_t�����[Ð��&    1����S[Ã���P�:Tt1�Ð�t& V��S�P��������x-�C(�K;K}!�S�4I���K����t�B�   ��[^�1�[^Ít& ��'    �P�:_t�   �f�������c�������Í�    ��'    WVS�Í@�C���������   �{�C)�9���   �C�7�Cu=��	~��jh�4	W�� ����t1������v����C,[^_����������������8$u����C붍v �G<_��<.���u<$u��	Nu��C0�   ��4	��)��C0������렍�    1�뙍�    ��    1�농�    ��    ��VS��u!�@�8 u1�[^Ít& ��'    �P�S���ht2��vuݍs���3����S�:_u˃����S�������    ��    �C�����C�8_u����C�   땍v ��  ��tZ�A��@��t:�8/u5�� �#��&    ��'    �8/u��t'�@����u���t����'    1�Í�    ��'    �@�ǀ     1����������������VS�ƉӃ���t3�;Jw��$�`%	��t& �S���������u�[��u؍t& ��'    1���[^Ð��&    �S���&�����t�8/u݃�[^Í�&    WVS�t$�|$�F�^�D9�wG�F��t[^_Í�    ��    �F��W�t$P�'� ����F�  ~[^_É���'    �V��u���u��v2���&    ��'    �9�w���S�6�cg ����t��^�w����   �݃��6�G �    �F    ���F    �F   �J����v ��'    UWVS�ƉӃ�(R�C� ����tx��   �,�(��    ��'    �σ�����   �>9눖  tE���   �uڈT$����  h�   V1�Ɔ�    ��  ����   �   �T$�f���[^_]Ð��&    UWVS�Ã�@Rh�4	�l$#U�~ �,$蓊 ������   ��   1��%�v ��'    �׃�����   �;9ƈ�  tU���   �L5 u؉D$�L$����  h�   1�Sƃ�    ��  ����   �   �D$�L$띐��&    ��<[^_]Ð��&    U��WVS�Ã�|�ɉU��M��w  ��  ����   �E�� ��K��  �$��&	�}�1��W�:'u4�R�r��r)����   ��u�}��W�
��u�zu	��;�O&  ��   =�   �   �P��   �(�E�ƃ  (�U��H���N�����   =�   ��  �P��   �)�E�ƃ  )�8<��!  ���Z!  �E��U��H�������t& �e�[^_]Ë}��W��  �   ��  �P�؉M�������tH�8/��  ��  �}����    ��    �@����t�8/u�� �}�u�@���|  ��t�E���  ��������������ǃ     �e�[^_]Ë}��u��؋O���L����غ�6	������O����4����]   ���x����#����}��u��؋O�������غ�4	�����O���������]   ���=���������E�1��P���)������M��&$  ��&    ��'    �8/�z  �P���o  �@����u�A�E��G��E�1��E���u��M��؋U���  �z���9u���  �E���   �6	�E��1��&    ��'    �у�����   ���6	��  �]  ���   �u҃���  �E�h�   Sƃ�    ��  ��   ���   1��E�롉غ�5	�����E��U��H�������������غ�6	�_����E��P�؃�������}   �������������   ��6	�}��1��&    ��'    ��������   ����6	��  ��  =�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢋�   ��6	�}��0��    ��'    ��������   ����6	��  �'  =�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢋�   �h6	�}��0��    ��'    ��������   ����6	��  ��  =�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢋�   �M6	�}��0��    ��'    ��������   ���W6	��  �  =�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢋E����p�E�h�4	P�ǉE��bx �����������!�%����t�M������  DWD� �����)��E�����   1��M��'���&    ��������   �9���  �����M�=�   �1uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢋�   ��5	�}��0��    ��'    ��������   ����5	��  ��  =�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢋E��P��   =�   �\  �H��   ���  �����}��u��؋O�������O�������������E��x�@�E���}���1��  ��3��  �M��U����\3  �M��U�����3  �����E��U��H���:3  ������   �6	�}��(��t& ��������   ���!6	��  �|  =�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢋E��6	�@���x��   �M��%f���������   ���6	��  �[  =�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢋�   �6	�}��0��    ��'    ��������   ���!6	��  ��  =�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢋E��H��t
�U��������E��@��������   ���   �(  �E��6	�E��/��    ��    �������   ���6	��  �2  ���   �u҃���  �E�h�   S�   ƃ�    ��  ��   ��1��E�롋E��H�p��t
�U����e����غ{   �����U��؉��M����}   �������<����E�f�x
 ��  �E��H�y�2	t�U��������    ���Y����E�f�x �  ��5	�����������ǃ     �������   �>6	�}��.�t& ��'    ��������   ���L6	��  �  =�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U��ǃ     �N����E��@�87������}���w�}���zc��  �}��?1�  �ֹ   �(6	�Hu	�9�   �U����%0  �E��   �+6	�@�P�E�������������8��  �   �ֿ(6	���  �E��U��@�H����/  �E��@�81������@�x������@�8>�x����)   �������g�����&    �E��@�89������P�::������@�}��   �E��B��E��B�}��E��G�.6	�0���  �غ56	�����E��x t�U������"/  �    ���6����}��M��؉�������E����������������.  ������    ��    ��  �}��U��E�    �E��E��}���  ��  �O�E����{����U���u�M��U�����  �E���  �Y����E���  �U��E�    ���E���  ��  ���}��U��E���  �G� ������  ���   �}��U��M����P�����wT�x��uG����  �8������L��|��x�y�x�y�x�y��  �L�U���  �@   � ��u��E��U��}��E��E��H�������M���  ���u�����t;�}������|�E��E��E��E���U����؃���  ��u�E���  �E��M����U�W�؃��q$  �������E� �<  �E��@��t
�E�@��  �M��U�����  �؃�����&  ��������E��U��H�������������غ35	�V����E��U��H�����������غ/5	�5����E��U��H�����������غ5	�����E��U��H���d����_����غ5	������E��U��H���C����>����غ�4	������E��U��H���"��������غ�4	�����}��u��؋O��������غ�4	�����O��������������غ�4	�v����E��U��H�������������غ�4	�U����E��U��H�����������غ~   ������E��U��H�����������E��U��H���o����j����E��x��   ���,	  �\6	�2����������������������   ���`6	��  ����=�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢋U��؃��������X����8/�3  ��  ���؋��  �U�������  ������<  �E���  ǃ      �E��E��}���<  �@t�0��u
�x�|  �U������P�����  <�x  �<   �������E��U��H���'�����  >�>  �>   ���^����E���  �E���<  ������E��x�p���������   ��+��    ��    ��������   �9���  �����=�   �u׃���  �U�h�   Sƃ�    ��  ��   ���   1��U�릋�   ��5	�}��$���������   ����5	��  ��  =�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢋E��}��H�������������t  ��4	���u����E��H�9E��  �U������������E��E��j  �x�p���������   ��!f���������   �9���  �q���=�   �u׃���  �U�h�   Sƃ�    ��  ��   ���   1��U�릋�  ǃ      �E��E��x��tW��  �M�1�1��E��E��M��E��M������E���  �x�H�@    �J����  ���t�����U�u�ǃ     �����E��E��@�B  �x�0���������   ��&��&    ��������   �9���  �a���=�   �u׃���  �U�h�   Sƃ�    ��  ��   ���   1��U�릋E�1��@�8��  ���#�$  �}�;�  ��$��  ��  �t& ��'    �E��}��E�    ��  �E��E���  �E��E��H�U��������E����T  �E�����  ������E���  �����غ�5	�����E��U��H���h����c����غp5	������E��U��H���G����B����غ`5	������E��U��H���&����!����غE5	�����E��U��H������� �����  1�������  ���^  ���v �J��u�J�	�q��w9��#	  ���u�1��������   ��5	�}��*��&    ��������   ����5	��  �2  =�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢉غ�5	������E��U��H���!�������ǃ     �����~������N�9>������غ(   �;����}��G�@�0�G�������&    �E��E��E��E�9��+��������O�U������������O�U������������M��q�M���Q�����  1��|>� ��)��h�����   ��-��&    ��'    ��������   �9���  �1���=�   �u׃���  �U�h�   Sƃ�    ��  ��   ���   1��U�릋U��O���4!  ������O�U��������������O�U����������   =�   ��  �P��   �)ƃ  )�����O�U��������������U��H���u����غ�6	�	����W�؃������}   �������K������U���4	�H���7�����   �.����������������������   ����4	��  t@=�   �u׃���  �U�h�   Sƃ�    ��  ��   ���   1��U�릋O�U������������O�U������������O�U������������E��U���   �H���u���9�   �i���9�   �]�������   �O����M��U�����  �����A���E�������*����a6	�"�v ��������   ���g6	��  t@=�   �u׃���  �U�h�   Sƃ�    ��  ��   ���   1��U�릍E���Wh�4	P�ǉE��d �����������!�%����t�������  DWD� ���   ����+}�tm�M�1��M���t& ��������   �9���  tD�M�=�   �1u׃���  �U�h�   Sƃ�    ��  ��   ���   1��U��=�   ��  �P��   �}ƃ  }�������   �6	�#��������   ���6	��  �����=�   �uӃ���  �U�h�   Sƃ�    ��  ��   ���   1��U�뢺.   �����������x�p���N�����   ��#�t& ��������   �9���  �!���=�   �u׃���  �U�h�   Sƃ�    ��  ��   ���   1��U�릋�  �E�������}��u�����  �؃柍O����  �O��������������������=�   ��	  �P��   � �E�ƃ   �p�������   ��5	�}��.����������������������   ����5	��  t@=�   �u׃���  �U�h�   Sƃ�    ��  ��   ���   1��U�릉}������G�   �"6	�0�E��u�� �u	����	  ��7�e
  �M��U��ؿ%6	�:  �u��   ���  �u���7	�   ��������   =�   ��	  �P�M���   �U��(��ƃ  (�S�����   =�   �D	  �P��   �)ƃ  )�)�����(  ��$  ���}�~+;�����}�1ɍW��t& �׃�;B��������9�u�;�,  �y	  �}�����  ����(  ���B����}�ta��4  ��8  ��    9��u��M��6	  ��|����M���E�;}��	  �u��0  ���A�F�2��	��u׋�|�����4  �    �P��1��������r����������    ��'    ��   =�   ��  �P�M���   �U��(����ƃ  (�K  ��   =�   �/  �P��   �)ƃ  )��������  �3 VS1���  ǃ       ��   �������E��U��H������������  ��t& �@���������8/������� �������@��������������&    ��'    �p�x�9�rB�/�������������������   =�   ��   �H��   ���  ��9���������)���~ƀ�_u��~_u��~Uu��F9ǉE�v�1����&    ��0���E�E�9��+  �E�� �HЀ�	vۍH�����  ��7�̓���  �U�h�   Sƃ�    ��  ��   ���   1��U��E���ǃ     �B�����4	�؉M�������M��A�P���c�����4	�������M��I�F�������  ƃ�    h�   S��  ��   ���   1��.�������  �U�h�   Sƃ�    ��  ��   ���   1��U��o�������  ƃ�    h�   S��  ��   ���   1��6�������  ƃ�    h�   S��  ��   ���   1��������  �}��U��E�    �E��E��}��⟉�  ��  �O�E��������E���  �E���������    ���6���������M��U��������������}��W�:���<�����<�  �E��U����H��������������$��'	�	���'���������	�������q����l   �������`����u   �������O����:6	��������>�����&    ��'    �H��  �E�    �E��E��ɉ�  �E��E���  �E��E����:������&    �H�����  ��W�����    ��� ��������    �������w����غ[   ������E��U��H�������]   ������������-   ��������_����:�O���v��c�����<����}��M��؉���  �غ<   �����u����F�H���6����غ�6	������F���H�������)   ���_����
�������  ƃ�    h�   S��  ��   ���   1�������E����E��O  ���X  �O�9E�@  ������>  ����������}��}���E������������P�  ���H�P�P��@�    �P�P��x��P�P���I�����v��E��}��U��H���4����?��   ��t9�}������|������t$�����u��غ    �M����O��U����  �ՋE���  ������p��4	�   ��o����E��U��H�������l8	���O��������غ[   ������E��U��@�H�������]   �������������E��}��E��E���  �E��U��H���X����?�(����E���  �����E��U��H���1����}� ��  ����������M��U����  �W���P��  h�   Sƃ�    ��  ��   ��1��Q����A�8)t
ǃ     �I�U�����  �����P��  h�   Sƃ�    ��  ��   ��1�����P��  h�   Sƃ�    ��  ��   ��1��F����}��M��؉��  �M�������  �M������n  �غ16	������M������V  �!����E��@�8�V����}��W�:)EǉE��B���P��  h�   Sƃ�    ��  ��   ��1�����P��  h�   Sƃ�    ��  ��   ��1��4����E��U��H����  �X6	���,�������1�1������_   �T����I������4  ǃ     �W����E��}��H�����u  �M�������  �4����B� <0��   <1�������	����������;}�v�<_u����   �z�����   �   ��u.ƃ�    P��  h�   S��  ��   ǃ       ����   ��u��P��   ���  �����-   ��������������	�������x������&    UWVS���9�w���*w;�͉׉��$��'	f���   =�   ��  �P��   � ��ƃ   �M�؃�[^_]�������&    ��   � 7	�&�v ��������   ���
7	��  ��  =�   �uӈT$��ƃ�    ��  h�   S��  ����   �   1��T$렍t& ��'    �I�d������&    ��   ��6	�&�v ��������   ����6	��  ��  =�   �uӈT$��ƃ�    ��  h�   S��  ����   �   1��T$렍t& ��'    ��   ��6	�&�v ��������   ����6	��  �  =�   �uӈT$��ƃ�    ��  h�   S��  ����   �   1��T$렍t& ��'    ��   ��6	�&�v ��������   ����6	��  ��   =�   �uӈT$��ƃ�    ��  h�   S��  ����   �   1��T$렍t& ��'    ��   ���   ��  �B��   � ƃ   =�   �/  �P��   �&ƃ  &�t& ��'    ��[^_]Ð��&    ��   ���   ��  �B��   � ƃ   ��6	�"�v ��������   ����6	��  t�=�   �u׈T$��ƃ�    ��  h�   S��  ����   �   1��T$������������������G�����   =�   �r  �P��   �*ƃ  *������    ��'    ��   �������t& ��   �+�����t& ��   ��6	�&�v ��������   ����6	��  �����=�   �uӈT$��ƃ�    ��  h�   S��  ����   �   1��T$렍t& ��'    ��   ��6	�&�v ��������   ����6	��  �=���=�   �uӈT$��ƃ�    ��  h�   S��  ����   �   1��T$렍t& ��'    ��  (t%��   =�   ��  �P��   � ƃ   �M�؉���6	�a�����   �,����'    ��������   ����6	��  �}���=�   �uӈT$��ƃ�    ��  h�   S��  ����   �   1��T$렍t& ��'    �M�؉��������   =�   ��   �P��   �)ƃ  )������v ��'    ��ƃ�    ��  h�   S��  ��   ���   1�������ƃ�    ��  h�   S��  ��   ���   1�� �����ƀ�    ��  h�   P��  ��   ���   1�������ƃ�    ��  h�   S��  ��   ���   1�������ƀ�    ��  h�   P��  ��   ���   1�������ƃ�    ��  h�   S��  ��   ���   1��������ƃ�    ��  h�   S��  ��   ���   1��_���f�UWVS�˃�<�ɉT$�l$Pty��  �ƅ�t�k��    ��'    ��  ��uT�S��uG�K��u�P��v6�S��)�C   ��  ��  t)��*tH��tg�T$���N�����  ���u���<[^_]Ã��3���T$���  ����  ��<[^_]Ã��3���T$����  ����  ��<[^_]Ë�  �T$��ǆ      �I�D����D$��  ��   uj��4	�\$�%��    ��������   ����4	��  tW=�   �] uփ�Ɔ�    ��  h�   V��  ��   ���   1��=�   tX�P��   �.Ɔ  .��\$�C�X���Eu�a��&    �[�����v�T$�ى��v�����  ��<[^_]Ã�Ɔ�    ��  h�   V��  ��   ���   1��y�����   ��4	�\$�������   ����4	��  t:=�   �] uփ�Ɔ�    ��  h�   V��  ��   ���   1�묋\$���C��Ph�4	�D$#P�L X�D$#P�X ������   tm1�\$����ȃ�����   �9Ո�  tD���   �\,u؉T$��Ɔ�    ��  h�   V��  ����   �   1��T$릋\$��4	�\$��ȃ�����   ����4	��  t;���   �] uՃ�Ɔ�    ��  h�   V��  ��   ���   1�뫋\$�,�����    ��    UW��VS�Éփ��D$0���G  ��&    �P����   � ��u���؉�j �L$@�-�����   ��=�   �9  �P��   � ƃ   ���   ��  �B��   �[ƃ  [���t�؉�������   =�   �%  �P��   �]ƃ  ]��[^_]É���'    �@�8*��  ��   �U6	�&��&    ��������   ���W6	��  tQ=�   �U uֈT$����  h�   Sƃ�    ��  ����   �   1��T$룍�&    ��'    �����j �L$@�������   �����   t�B��   �)ƃ  )��������  ƃ�    h�   S��  ��   ���   1�뻐�t& ����  ƃ�    h�   S��  ��   ���   1�������&    ��'    ��ƃ�    ��  h�   S��  �[ƃ  [�����   ǃ      ���=����   �M���f���   �������t& �����j �L$@�������   �����������  ƃ�    h�   S��  ��   ���   1�������&    ��'    UW��VS�׉Ã��t$0����   �F����   ��   �\$�-�����������������W  � ����   �H����   �H�	����wމ�����1 ��tǋ\$��  < �-  ��   ���   �V  �B=�   ��   � ƃ   �  ��ƃ�    ��  h�   S��  ��   ���   1���   ��\$��  ��ǃ      ����D$j ��������   �����   �	  �B��   �(ƃ  (�M ��t�؉�������   =�   �.  �P����   �)ƃ  )j�؉�������D$����  ��[^_]Ð�t& �\$��  �����(�������   =�   ������P��   �(����  ƃ  (��ǃ      ���D$j ��������   ��=�   ��   �P���   ��   �)ƃ  )�������ƃ�    ��  h�   S��  �(ƃ  (���M ��   ǃ      ��������   ������t& ��'    ��ƃ�    ��  h�   S��  ��   ���   1�������ƃ�    ��  h�   S��  ��   ���   1��%�����ƃ�    ��  h�   S��  ��   ���   1��{����v ��'    WV��S�É΃���<  ��t��  �D$�T$�T$��  ��9t+�����r�����<  ��t
�D$��  ��[^_Í�&    �I�؉��D�����<  ��t
�D$��  ��  <��   ��   =�   tf�P��   �<��ƃ  <��H���������  >��   ��   =�   tj�P��   �>ƃ  >��[^_�������������������  ƃ�    h�   S��  ��   ���   1��k�����&    ��'    ����  ƃ�    h�   S��  ��   ���   1��g�����&    ��'    ��   ���   tI�B��   � ƃ   ���������'    ��   ���   tH�B��   � ƃ   ���������  ƃ�    h�   S��  ��   ���   1�닃���  ƃ�    h�   S��  ��   ���   1�댍t& ��'    �91t�f�����    WVS���Q�z�r��tm�����   ����������   �9���  tE=�   �uۈT$��ƃ�    ��  h�   S��  ����   �   1��T$먍v ��[^_É���'    UW��VS����T$��0���������Ɖ����ui��td��   �T$��=�   tq�p��   �(��ƃ  (�v�����   =�   ��   �P��   �)ƃ  )��[^_]É���'    �T$����[^_]�.�����&    ��'    �L$�T$��ƃ�    ��  �   h�   S��  ����   1��L$�T$�P�����&    ��'    ��ƃ�    ��  h�   S��  ��   ���   1��<�����&    ��'    �H�9Lt1�Ð�t& UWVS�Y�ƃ��X�Q��_����Z��   ����   ���/I  ����tr�8'��   �V�;   �<n��   <E��   ��tJ�Z���    ��    ����t2�^�<Eu��)щ��4��������P��蕷���^�����EtG��1�[^_]Í�    ��'    ��u<1���Zuك�1҉��^�h  �^���Eučt& ��'    ���^��[^_]�f��Y�^�Q븍t& �Jf�< �N�B���.����t& ��'    �@�P�������@)F0�����1��5���UWVS��<�p,�H�t$�1�V�����  �Q�ŉP�A<E�Z  �D$,    �\$,�Y��&    ��'    ��I<�%  �����������\  ���/   ��j �c���������>  �U�X�<E�e  <L��   ~�<X��   �E4�z�E4   �}�$�B<L�T  <T�l  <s��  <f��  �HЀ�	��   <o��   <t���U  �zl�S  ����[  ���D$�@  �D$� ��1��   ��2�h  ��3�  �E�8_�c  ���E   �E���q  �S  ��    ��    ���)����������f����F  �������f��zn�s������U���]  ���U��   �:I���  �$�E4�:Et1���<[^_]Í�&    ��'    ���U�y�����t& �D$�   �@�x�0�W�U0�t$��7	��!  �@����  ��  ����  ��u(�t$�.6	�   ��  �D$�8n�  ��t& �U1��S�����    �B<r�M  <p���������U�/k  �����I   j ��   ��&    ��'    �zp�S����B�E�zT�3  ���U1ҋE;E}��u�@���E����t	�   �Q�U����f��D$���U�E,�D$,��<[^_]Í�&    ���y����U�����������������������ɹ���U���l�����������������1�����  �G�E   �E���T  ����0   P���R����U�����"�����t& �D$�@���   ~.�D$    �k�����D$���5������   P�L$뭍�    ���x������4   j �L$돋D$�@� �xc��  ���i  �D$�t$�(6	�   ��d  �t$�7	�   �t�t$�7	�   ��u  ���eZ  �ƋE�8I�Q  ���7   ��V�L$ �c����L$�$�6   ��������/   ��Mj 1��<���Z� ������E���	i  ���5   P�L$��������U�:C  �ǉ���Y  �ƋE�8I�+  ��V���   �������̷������������L����D$� <mt<pu��|$:Gu��E�8_�r������h  �����7   P��菱���L$�$�5   �%����@<at<w������_   ���R  �D$���B  �U�D$�<E��  1�<p�$  <i�����zl��������U�E   �  ��1�P�0   �������������:   ��Q�L$�����L$ �$�9   ���ٰ���L$�$�8   �o��������������   P��诰���$��������A  ���5   P�L$�5������A  �}�������U�<L��  <T��  <s��  <f�c  �HЀ�	��  <o��  <t��t<iu
�zl�W  ���GV  ���D$��  �D$� ��1��  ��2��
  ��3��  �E�8_��  ����f  ���5   P�L$���ӯ���D$ �E�����L��  ��T�L
  ��s�  ��f�L  �JЀ�	�D  ��o�+  ��t��t��iu
�xl�Q  ���U  ���D$�R  �D$� ��1��  ��2��  ��3�1  �E�8_��  ���f  ���5   P�L$�������D$�E�����L��	  ��T�  ��s�]  ��f��  �JЀ�	��  ��o��  ��t��t��iu
�xl�4  ����T  ���D$��  � ��1�;  ��2�  ��3�c  �E�8_��  ���[e  ��P�L$$�5   ���g��������]�����    ��'    �E   ���4  �������� �P���v��c<�R������P?  �D$�M����U�<L�  <T�q  <s�M  <f��  �HЀ�	��   <o��   <t��t<iu
�zl�h  ����S  ���D$��  � ��1��
  ��2�y  ��3�d  �E�8_�A  ���ed  ��P�L$�5   ���q��������������&    ��1ɉU�S����zn��������U���U  ������  �E�8I��������?�������   P���������������xn�;������E����T  ����������E�8I�������L$��������   P�L$$��跬�����������zn�u����B�E���vT  �D$���E��������I��������������   P�L$ �����xn��������E���+T  �D$���E��+�����I�"������I������   P�L$������zi���������U�E   ��  ��������zp������B�E�zT��
  �B1ɉE�U;U��  �}�4R���U�<����|$������|$�   �O�������P��r��  ��p��������E���Sb  �����I   j ���`��������V����xp������P�U�xT��
  ��1ɉE�U;U�  �}�4R���U�<����|$������|$�   �O�������xp�0����P�U�xT��   ��1҉E�E1�;E������M�4@���E����������   �Q�����P��r�V  ��p�������E���`a  �����I   j �M����B<r�3  <p�-����B�E���.a  �����I   j �c������&��������U���1��$����E��D$    �K����E��D$    ������zp�,����B�E�zT��  ��1��U�U;U��  k��u���U΅��C����   �F�5����B<r��  <p���������U�k`  �����I   j ���x��������������&    ��'    �D$�@�������
  1҃���  ���%����ֿ.6	�   ��-  �:n�����B<at<w������_   ����  �Ɖ��$:  �ǋE���E��
  ��p��
  ��i��
  �xl��
  ���_  �����:   P��讨����$�9   ��蝨���L$�$�8   �j����D$��7	�@��D$�@�֍H�M0�   ���������8��  �D$�@���d  ��������'������4   j �L$����1�����  �E�E   ����  ����0   P��������$�����������������D$�E�����1����  ����U�E   �  ����0   P��������ԭ���D$�E�������D$�@��������   1҃��d  ���@����ֿ.6	�   ��A
  1ɀ:n�L����B<at<w�<����_   ���   �Ɖ��W8  �ǋE���E�?
  1ɀ�p�
  ��i�����xl���������]  �����:   P���ߦ����$�9   ���Φ���L$$�$�8   ��軦�������������~������4   ��j �L$$蔦����������1�����  �E�E   ���`  ����P�T����D$��7	�@��D$�@�֍H�M0�   ���������8��		  �D$�@���  �h�����������D$�@� �xc��	  ��T$��\  �T$�D$�(6	�ֹ   ���	  �7	�ֹ   �tPPh7	R�:: ������	  ���M  �ƋE�8I��  ���7   ��V�L$(腥���L$$�$�6   ���r��������h�����葫���D$�E��D������������D������-������X���1������D$�@���/����
  1҃��0  ��������ֿ.6	�   ��b  �:n������B<at<w������_   ���  �Ɖ���5  �ǋE���E�}  ��p�W  ��i�A  �xl�%  ���m[  �����:   P���{�����$�9   ���j����L$�$�8   �����D$��7	�@��D$�@�֍H�M0�   ���������8���
  �D$�@���W  ���������������4   j �L$�����������D$�E�������D$�@� �xc��  ��T$�Z  �T$�D$�(6	�ֹ   ���  �7	�ֹ   �tVVh7	R�8 ������  ���SK  �ƋE�8I��  ���7   ��V�L$ �Q����L$�$�6   �f������E���c4  �Ɖ��
K  �ǋE�8I�J  ��W��   ������<mt<p�{���:B�r����E�8_��  ����Y  �����7   P���Ϣ���$�P�����&    �D$�   �@�x�0�W�U0�t$��7	���  �@���  ��  ���|  ���@���WWh.6	�t$ ��6 �����  �D$�8n�����@<at<w�����_   ��� 	  �ǉ��W3  �ƋE���E��  ��p��  ��i������xl���������X  ����:   P���������$�9   ���С���L$�$�8   ��轡�������<����v �D$�@� �xc��  ��T$�rX  �T$�D$�(6	�ֹ   ���  �7	�ֹ   �tQQh7	R��5 �����w  ���'I  �ƋE�8I�w  ���7   ��V�L$$�%����L$�$�6   �����������������E�-���������v ��'    ���������k����<mt<p�����:B������E�8_�P  ���W  �����7   P��襠���L$�$�5   �r����t& ��蹦�����������k��������E�9����Z������&    1����"  ����U�E   �4  ����0   P���2������������D$�@��������a  ���D$    ������D$�@� �xc��  ����V  ��PPh(6	�t$ �V4 �����K  PPh7	�|$ W�:4 ����tPPh7	W�&4 �����k  ���sG  �ǋE�8Iu�����������   P���p������ǃ���7   W���Y����L$�$�6   ���F��������������    ��    �B�E���S0  �ǉ���F  �ƋE�8I��  ��V���   �"������E���0  �ǉ���F  �ƋE�8I�p  ��V���   ���ƞ�����������<mt<p�����:B������E�8_�r  ���qU  �����7   P�������L$�$�5   �������E�-����xi�%������E   �E���7  �O������E1��B����i   �D$    �N����D$    �����xiu����E   �E����  �9������E1��,���� �H���v��c<������T$��.  �T$�D$�������T  ���K��������������   P��藝��������������fT  �Ɖ��]T  �ǉ��TT  ������i   �D$    ������D$    �����xiu����E   �E���(  �������E1��������O.  ��P��������S  �Ɖ���S  �ǉ���S  �����xi��������E   �E����  ��������E1���������E   �E���  �8�������-  �U�����������������   P��艜�����������E   ���c  ������� �P���v��c<�h������-  ���c������q-  ���5   P�L$�������S  �������E   ���  ���u���� �H���v��c<�������T$�-  �T$�D$��������R  ���9���������������   P��蹛���$�������u������4   ��j �L$蔛�����������D$� <mt<p������|$:G������E�8_t?���;R  �����7   P���I����$��������R  �ǉ��R  �Ɖ��R  �0������E�������A,  ��P�����E   ����  ����������Q  �Ɖ���Q  �ǉ��Q  �������Q  �������E   ���  ���}���� �H���v��c<������T$��+  �T$�D$�����<i������������+  ���R������E   �E���K  �'������E��������E   �E���)  �������]+  �U����������E   �E���  �%�������U�/+  �ǉ���A  �ƋE�8ItM��V���   ���ڙ�������Y�������*  ���B��������������   P��詙�������f�������������   P��膙���$뙉��*  ���5   P�L$��������������   P���O����$�s������`�������   P���.����$�������E�-����t& ��'    UW��VS��<�X�D$,�T$�D$,    8�D$�w  �ڍ�    �]4�E4   �<L��  <T�  <s�  <f�S  �HЀ�	��   <o�   <t����  �zl�
  ���>  ���D$��  � ��1��  ��2�S  ��3�z  �E�8_��  ���'O  ��P�L$$�5   ���3��������i  ����'    �znu����U����?  ���%  �U���:I��  �]4���.   ��j �����|$�������   �U���D$�D$8������ӋD$,���]��<[^_]Í�&    �B<r��  <p��������U�_N  �����I   j ���l��������   f��zp������B�E�zT�6  ���/�����tZ�U;U}R�M�4R���U����t?�   �A������D$�@���������  ���!  ����  ���&    �]41���<[^_]Ív ����������&    �ɉ]4������֍v ���ٜ�����名t& �D$��7	�@��D$�@�֍H�M0�   ���������8��Z  �D$�@����  �T  ���}  ���b����.6	�ֹ   ���  �:n�E����B<at<w�5����_   ��������Ɖ��0'  �U���<E��  <p��  <i� ����zl��������L  �����:   P��轕����$�9   ��謕���L$$�$�8   ��處�������������������������1����v  ����U�E   �T�������0   P���R��������������&    �D$���U������   P�L$$���!��������W�����&    ��1��U������v ���������4   ��j �L$$����������������'    1ҋD$�@� �xc��  ��T$�K  �T$�D$�(6	�ֹ   ���  �7	�ֹ   �td�7	�ֹ   �tT���MK  �ƍt& ��'    ���7   ��V�L$(�L����L$$�$�6   ���9��������o���������������������;  �ƋE�8Iu����(�������   P������������������������������U�%  �Ɖ��;  �U�ǀ:I�*  ��P��   ��誓������������<mt<p�C���:B�:����E�8_�l  ���UJ  �����7   P���c����$�����t& ��'    1ҿ.6	�   ����������J  �Ɖ��
J  �ǉ��J  �M�����    ��    ���9$  ��P�������)$  �U���y������������������E   ����������m�����    ��'    � �H���v��c<�������T$��#  �T$�D$����������������   P���y����$�������.   1ɉ]j ���[���Z�z������E   �E���3����������1��U�b����zi�G�������U�E   �����A������E����<i�i����n������&    UWVS�Ã��@�8_t/���h����ƅ��n  �S1��:_��   ��[^_]Ð��&    �p�k4�C4   �s�P��L��  ��T��  ��s��   ��f�  �JЀ�	��  ��o��  ��t���/  �xl��   1����#  ���E   �؉s�!��������0   P�����������  ��t& ���؉S�3"  ����-   P����������[^_]Í�    �P��r��  ��p�-  ����6  ���$��  � ��1��  ��2��  ��3�{  �S1��<_�  <L�7  <T�=  <s�*  <f�k  �HЀ�	�`  <o�H  <t��t<iu
�zl��  ���[6  ������
  � ��1�  ��2�9  ��3��
  �C�8_�  ����F  ��P���5   ��������������  ���7   ��Q�ҏ���$�L$�5   ��迏�������5���&    �xn��������C���y7  �����o  �C�8I�3  �k4�����t& ��'    �xp������P�S�xT�  ��1҉C�C;C�"  �K�4@���C�4���t��   �V롍t& �$�@���g  ��  ���D$    �L  ����   �t$�.6	�   ��5  �D$�8n��   �@<at<w��   �_   �������ǉ���  �ƋC���E��  ��p� 	  ��iuj�xlud���]E  �����:   ��Q���i������$�9   ���X����L$�$�8   ���E��������������$����������������'    1���������'    �������������f����)������o���f��$�   �@�x�0�W�S0�t$��7	���  �@���  ��  ��������$�@� �xc�  �C���L�q  ��T�x  ��s�1  ��f�  �JЀ�	��  ��o��  ��t��t��iu
�xl��  ���_3  �����  � ��1�.  ��2�   ��3��  �C�8_��  ����C  ��P��5   �������D$���t$�(6	�   ��  �t$�7	�   �t�t$�7	�   ��V  ���4  �ƋC�8I��  ���7   ��V�L$腌���L$�$�6   ���r���������������&    1���������'    ���i�������   P���7�������������    ��'    ����������4   ��j �L$���������v������C���  �Ɖ���3  �ǋC�8I�k  ��W��   ���Ë�������6����D$� <mtX<ptT�S1���������C���pB  �����I   j ���}���������������؉S�E   �Q�������Q�����|$:Gu��S�   �<_��������S�f����Y  ��P�Q������I  �s��������zn��������S����2  ���������C�8I������؉L$��������   P�L$���Ê������������E   �������������C���L��  ��T�  ��s��  ��f�H  �JЀ�	��  ��o��  ��t��t��iu
�xl�>  ���i0  �����	  � ��1��  ��2��  ��3��  �C�8_�j  ����@  ��P��5   ����������ǋC���L��  ��T��  ��s�c  ��f�  �JЀ�	�V  ��o�=  ��t��t��iu
�xl�Z  ���/  ������	  � ��1�>  ��2��  ��3��	  �C�8_�]  ���A@  ��P��5   ���O������ƋC���L��
  ��T��  ��s�u  ��f�  �QЀ�	��  ��o��  ��t��t��iu
�xl�  ���/  ���D$�%	  � ��1��
  ��2�n  ��3�	  �C�8_�u  ���?  ��P�L$�5   ��蝈�����������v � �P���v��c<��������  �D$�~��������������   P���Q����$�x����B<r��  <p��������؉S�?  �����I   j �����������!����t& ��'    �zp������B�C�zT�`  ��1��S�S1�;S�����k�K���S��������   �A������xn�^������C���w/  ���D$�k  �C�8I��������������   P�L$���d����D$���l������1>  �������P��r��
  ��p��������C���>  �����I   j �������D$���������&    ��1ɉC�x����xp������P�S�xT��  ���C1��S;S��  k�K���S�ɉL$������   �A��������������   P��膆������������xn��������C���E.  ���������C�8I�������h�������   P���6�������������xn�.������C����-  ����������C�8I������؉L$�������   P�L$������������[����xn�|������C���-  ������  �C�8I�����������������   P��萅�������������o����������1������xi�E������E   �C���C�������������������T������g������F������������O����D$    �'����G��@QQh�7	��C0R�T$�u �����T$�]  �G�@����  ��  ���   ���H���PPh.6	R�T$�. �����T$��  �:n�����B<at<w�����_   ���i����D$���  �D$�C���E��  1ɀ�p��  ��i�]����xl�S������;  ���:   P�L$���"����L$�$�9   ���������$�8   ������������
����P��r��  ��p��������C���:  �����I   j ��较�����������P��r�0  ��p��������C���q:  �����I   j ���~�������������P��r��  ��p��������C���1:  �����I   j ���>�������������xp������P�S�xT��  ���C1��S;S��  k�{���S��������   �G������G���������  1҃�� ����G� �xc��  �؉T$�9  �T$�D$PPh(6	R�T$� �����T$�C  PPh7	R�T$�� ����tPPh7	�T$R�� ������  ���**  ���C�8I�.  ���7   ��Q�L$�(������$�6   �����������#����xp�����P�S�xT�'  ���C1��S1�;S�b���k�K���S���N����   �A�@����xp�����P�S�xT��  ���C1��S1�;S�A���k�s���S���-����   �F����1�����  �C�E   ���?��������0   P���=��������I���������������1��$�����������D$� ������5����D$�����F�8�@��C0PPh�7	W�b ������  �F�@���:	  �D  ����  �������PPh.6	W�# ������
  �?n�n����G<at<w�^����_   ���b����D$���  �ǋC���E�!  ��p��  ��i�$����xl�������7  �����:   P���!����L$�$�9   ��������$�8   �������D$���������s��������4   j �����������������赅���������1��:�����螅��������1��T���1���t	����  �ƃC�E   ���o�������0   P���m���D$���u������؉S�  �ǉ��+'  ���C�8I�
  ��Q���   ���+�������7����F���	�����  1����L����F� �xc�9	  ����5  �D$PPh(6	W�^ ������  QQh7	W�F ����tRRh7	W�2 ������  ���&  �ǋC�8I��  ���7   ��W�L$�}~����$�6   ���l~���D$���t������������������������������<mt<p�-���:B�$����C�8_�  ����4  �����7   P���~���$������������������D$�@��@��C0PPh�7	R�T$�O �����T$�  �D$�@�@����  ��   ���[  �������PPh.6	R�T$� �����T$��  �:n������B<at<w������_   ���?����D$���t  �D$�C���E��  1ɀ�p��  ��i������xl���������3  ���:   P�L$����|���L$�$�9   ����|���L$�$�8   ����|�������M������������4   ��j �L$�|�������&������C����  �ǉ��k$  �ƋC�8I�Q  ��V���   ���k|���D$���s����D$�@�������~�1҃�������D$�@� �xc��  �؉T$�3  �T$�D$PPh(6	R�T$� �����T$�+  QQh7	R�T$�l ����tRRh7	�T$R�T ������  ���#  ���C�8I�5  ���7   ��Q�L$�{���L$�$�6   ���{������������諁�����|�����蝁����������F�8�@��C0PPh�7	W�� ������  �F�@����  ��   ���  �������PPh.6	W� �����l  �?n������G<at<w������_   ��������D$���  �ǋC���E��  ��p�{  ��i������xl��  ���}1  �����:   P���z���L$�$�9   ���xz����$�8   ���gz�������e������2�������4   j ���Bz�������@����F������~�1���������F� �xc�_  ����0  �D$PPh(6	W�y �����)  PPh7	W�a ����tPPh7	W�M �����6  ���!  �ǋC�8I�
	  ���7   ��W�L$�y����$�6   ���y�������������U�������4   j ���by���D$���j���������������1����I	  �C�E   ����������0   P���y�����������1����X  �C�E   �����������0   P����x�����������1Ʉ��S  �C�E   �؉L$�������0   P�L$���x�������%����F���,�����   1҃���  �������PPh.6	R�T$�� �����T$�5  �:n������B<at<w������_   ���%����D$���Z	  �D$�C���E�^  ��p�3  ��i�`����xl�  ����.  ���:   P�L$����w���L$�$�9   ����w����$�8   ���w�������h�������������4   j ���w�������C����<mt<p�r���:G�i����C�8_��  ���B.  �����7   P���Pw���$�G����F��@QQh�7	��C0R�T$� �����T$��  �F�@���
  �S������y����F� �xc��  �؉T$��-  �T$�D$PPh(6	R�T$�J �����T$�T  PPh7	R�T$�* ����tPPh7	�T$R� ������  ���_  ���C�8I�  ���7   ��Q�L$�]v����$�6   ���Lv������������E   ���&�������������C���R  �ǉ���  �ƋC�8I�&  ��V���   ����u������������E   ����������K������,  �D$���,  �ǉ��,  ����� �P���v��c<���������  �D$�������  ���)������  ��P�{������C���  �Ɖ��B  ���C�8I�:  ��Q��   ���Bu��������������a  ��P�'����؉L$�=������   P�L$���	u���$������<mt<p�����:B������C�8_�  ���+  �����7   P����t���$�_����<mt<p�����:B������C�8_�  ���q+  �����7   P���t���$��������C���  �D$���?  ���C�8I�M  ��Q�L$�   ���=t�����������<mt<p����:G�����C�8_t����*  �����7   P����s���$������ �H���v��c<�$����؉T$�  �T$�D$�������*  �D$���*  �D$���*  �l������{*  ���X������C�s������C������؉L$蓼�����   P�L$���_s����������� �H���v��c<�����؉T$�d  �T$�D$������� *  ���f������C�����؉L$�#������   P�L$����r���������������������   P����r���$�����E   ������������� �P���v��c<���������  �D$�������d)  ����������E   �C���[����a������  ��P������xi�,������E   �C���*����������C1��������i������P����؉L$�/������   P�L$����q���$�������E   �C���������������C�i������(  �D$���(  �D$���(  ��������  ��P������xi��������E   �C���s����H������C1��;����xi��������E   �C���E����D������C1��7������E   �C���!����{������E�������   P���q���$�������E   �C����������������������   P����p�������@����E   ���������������'  ����������  ��������軹�������   P���p��������������  ���������C�Z����E   ���J����������� �H���v��c<�P����؉T$�b  �T$�D$�K�������&  �D$����&  �D$����&  ��������&  ���������  �������i   1�������xi�p   u���E   �C��������������C1��������E   �C�������������n&  �D$���c&  �ǉ��Z&  ��������   ��P�Z����؉L$�z������   P�L$���Fo������������xit1��v������C1��������E   �C��� ����n����i   �Ή؉L$�������   P�L$����n���$������    ��'    UWVS�Ã�,�h�E <V��<r������  <K�  �PЀ�J��   ���$�|(	�{4�C4   �E<L�0  <T�  <s�6
  <f��
  �PЀ�	��	  <o��	  <t��t<iu
�}l��  ���N  ������  � ��1�  ��2��  ��3��  �C�8_��  ����$  ��P��5   ����m���������{4�A   j ����m���D$,����t�S�: t�J�K�:E��   ��&    1���,[^_]Í�    �T$1ɉ��cn������t݋C�8F��tC�������tȋ8�O��v>�T$��t��C ;C$}��K�����C �D$��,[^_]Í�    ��  �뻍�&    �L$�x�H��T$�>뮍�    ��    �M�؉K�s�������(   j ����l���D$,������'    ���(����S ;S$�����K�����D$�S ��,[^_]Ít& ���y  �D$�Ív �U�S�E<_��  ��0<	��  �E�ƉC���>�OЀ�	v�)։؉���l������t�S�:_�Q  1���   ����'    �M�؉K�S��������%   j ���l���D$,���4����t& ���  �D$� ����M�؉K���������&   j ����k���D$,��������t& �E�C�} �����E�C�E��F<0��������$��)	��M�؉K���������9������������*�������+   P���Xk�����D$�|�����    ��    �M�؉K�c��������$   j ��� k���D$,���D����t& �M�؉K�3��������"   j ����j���D$,�������t& �M�؉K���������#   j ����j���D$,��������t& �E�PЀ�	v<_t��A<��  1҉���l���S�D$�:I�������蕳�����   P�L$,���aj���D$,��������t& �M�؉K�q���D$�Ɖ��f��������!   V���$j���D$,���H������&    �S;S�������4� 2	��  �C�<R���S������  �M� '   �p�VS0�K�'�����t& ����o���s�D$�>I������S8����  ��������S ;S$������K�����؉S 藲��������S;S�f  �C�R���S�����O  � '   �@l4	�C0�����S;S�-  �C�R���S�����  � '   �@D4	�C0�b����S;S��  �C�R���S������  � '   �@4	�C0	�)����S;S��  �C�R���S������  � '   �@04	�C0
������������-����S;S�v  �C�R���S�����_  � '   �@X4	�C0�������r��������I   j ���/h���D$,���S����S;S�  �C�R���S�����   � '   �@�4	�C0�L����S;S��   �C�R���S������   � '   �@4	�C0	�����   �7	���0h��������C;C��  �S�4@���C���T$�,   �E��0<	���Ȅ�f�Jt�C�gl���t$���|����F�D$�@��������C�Bl���C1Ҁ8 t�P�S1Ҁ8s�D$f�P
�o�����    ��'    �D$    �   1����؉S���������*   P����f�����s������  ���D$�����8������	����s4�C4   �E<L�S  <T��  <s�)  <f�i  �PЀ�	��   <o��   <t��t<iu
�}l��  ���i  �����]  � ��1��  ��2��  ��3�@  �C�8_�
  ����  ��P���5   ����e�����ǅ��s4�����1�������    �C(�k�{ �D$�C0�D$�������K�9I�R  �D$�s�k�{ �C(�D$�C0�D$������        �}n�3����M�K���V  ������  �S�:I�'  �s4�����E<r�<  <p������M�؉K�  �����I   j ���$e�������"����v ��'    �}p������E�C�}T�  �M1��K�S;S�   k�{���S����   �G�   �S�]����}n�~����M�K���  ���^  �S���:I������D$��襭�����   P�L$���qd�����������L$��������S ;S$������s�����S ���������������8����E<r��  <p������M�؉K��  �����I   j ����c��������������i����������s41��������j����������}p������E�C�}T�^  �M1҉K�K;K�\  k�C���K1Ʌ�������    �P�������G���T�����  1���@  ���n���QQh.6	U���  �����*  �} n�L����E<at<w�<����_   �������D$���7����ŋC���E��  ��p�m  ��i�����xl��������  ����:   P����b���L$�$�9   ���b�����$�8   ���b����������1����E  �C�E   ���i��������0   P���gb�������e����G�(�@��C0PPh�7	U���  �����I  �G�@���X  ��   ��������G� �xc�M  ����  �D$PPh(6	U�s�  �����P  PPh7	U�[�  ����tPPh7	U�G�  ������  ���	  �ŋC�8I��  ���7   ��U�L$�a�����$�6   ���a����������������������4   j ���\a�������Z������;g�����������1��\������R��������   P��� a�����������F�(�@��C0PPh�7	U�|�  ������  �F�@����  �b  ����  ��u�RRh.6	U�A�  �����z  �} n�k����E<at<w�[����_   �������D$�������ŋC���E��  ��p��  ��i�!����xl�������0  ����:   P���>`���L$�$�9   ���+`����$�8   ���`�������3����M�؉K�3����ǉ���  �ŋC�8I�  ��U���   ����_������������E <mt<p�����:E������C�8_��  ���  �����7   P���_���$����1����p  �C�E   ���`�������0   P���^_�������w������}e�����i�������������[����F���1�����   1���I����F� �xc�X  ����  �D$PPh(6	U�u�  ������  PPh7	U�]�  ����tQQh7	U�I�  �����/  ���  �ŋC�8I��  ���7   ��U�L$�^����$�6   ���^�������������1�������4   j ���^^�������w����E <mt<p�I���:E�@����C�8_�D  ���  �����7   P���^���$��������  �D$����  �ŉ���  ������������P����������������   P����]���$������ �H���v��c<�������������D$�����E   ���{�����������M�؉K�����Ɖ��N  �ŋC�8I��  ��U��   ���N]�������g������m������������_�����P�6�������  ���r����E   ����������]�������������   P����\�������:����xi��������E   �C�������q������C1��d���� �H���v��c<�������������D$�������g  ��������xi��������E   �C���T����������C1��������E   �C���0����G������  �D$���	  �ŉ��   ��������C��������9������������E   �C���������������C����������������   P����[�������������֤������   P���[���$�@�����    ��    UWVS���h�D$    �U ��E�������ut��.to�Ít$�L��&    ��'    �����.   j ���=[�������t=�k�p�U ��E���҉������u7��.t2��Ot��Ru�}Et"���+�����u�1���[^_]Í�    ��'    �D$��t�P��u܋P�:'uԋR�z	uˋR)S0�@    뼐VS�Ã��@�8Jt11���u1��������t@����)   P���~Z������[^Ð�t& ���C����������u�    ��'    1��э�    ��    �P�:Ft1�Ð�t& S�J���H�zYu���P�ú   �^������\���S�:Et��1�[Í�    ���S��[Ð�t& UWVS���D$�@�8 ��   �|$�P�W�x �8��   �\$�P�S�@����v�D$��   ��0<	wU���G`���K;K��   �S�4I�����K����   ����   �L$�B���2   ��0�J�z�t& �D$ 1��=   1҉\$���    ��    ��8�~E�D$;T$tD�D$��)Љ������Љ����� .	�� .	�8�u��N8L$t{:L$��P;T$u�1���[^_]�f��D$ 뀀|$v�u�����c�l����S41��s8�����C8���������s8��j �غ3   �xX������[^_]Í�    ��'    �D$�P;P}��ǋ@�R���W�����o���� 1   �h��[^_]Ív ��'    UWVS�Ã��@��JЀ�	��   �J�����   �J�����  ��L��  ��U�  �P��l��   ��t��  �P1�S�H��tuc���C���]������   �S;S})�K�4R���S�,���t�E�C ;C$�E F   �  �S1��
��t& ���^���S���
��B��t
��[^_]�f����؉S��]������J   P���!W���S���ŀ:Bt���f����)�������t	�81�:  �S�
�f��P1�S�H��lu����C���B����S�����
�q�����E�h������؉S�\�����6����S;S�*����K�4R���S�,��������}�E�C ;C$�E D   ������S�,����C �]�����&    �{,���|$t�7����   ����  ��C�Y  ��DuT�p�VЀ�wH���$�l*	��&    ��'    ���C���\������t���v\�����������&    ��'    ��1�[^_]Í�    �P�7	�   �BC0�2���C0���������V\������5   P���U���S�Ń��
�#����t& �WS0���C��   ��D�1�����1�������   �s;s�P�S��   �{�,v���s�,�����   �t$����   �M�t$�E    �u�H�������&    �   뢹   뛹   딹   덍t& �p�Vπ���������$��*	�   �s;s�P�S}c�k�<v���s�l� ��tO�|$��tG�M�t$�E    �u�H������    ��'    �   먹   롹   뚹   듍t& �H1�������t$�VS0������v UWVS�ƃ�,�@���S��  ~f��UtA��Z�(  ��1҉F���  �V�À:E�+  1ۃ�,��[^_]����������������������Ã�,��[^_]Í�    ��'    ��N��   ���T$�   �F���aT������t�1҉�1��pU���V�D$���    ��t|��D��  �C�<	��  �C�<�}  ��C����U����i  ��L�`  ��S�'  ��I��  ��T�E  ��E�g  ��Mu��t�B�F�Z��u��v �E     1������f��������V�À:I������������F ;F$������V�����F ��贛������P�8��    ��    �xttJ1҉���T���ǋF���8I��������z�������P�   ���HR������������&    ��'    ���F�������   �ú(7	���R�������   S����Q���ǋF�F0�����8I�0����������F ;F$������V�<����F �a���f�����������   �   ����P���Q�����ǀ�St(�V�:EtM��������F ;F$������V�<����F �V�����f��B���<T��u3�~�����u��V�ǀ:Eu��E   �������    ��뒍�    ��    ������ˉ���'    ���(������!����   �K�����&    �   ���DS�����+����V����o���������������������V���f����t& �B�F�B<s��   <dtK���s�������t� ��Dt��F��   ��    ��'    ��W�ى�   �^P�����Ã�,��[^_]Ã����V�2V�������]�������������t� ��Dt��Fu+�F1�;F}��N�<@���F�<���t��E   �o�W넉��T$�yV�����T$u�1��������cV�����[���1�����������V�GV����������   �7	���.P����P�)������} ������L$��t�D$�L$�A�F�8E��������\$�F������    ��    UWVS�Ã��@���T��   ��G��   �؉���������t
��t�CtI�C� <E�����ub��t^������   ��   ������   �R��u���   �v �v��P��v��u�V�����w��R�����v�V����[^_]Í�    �K0�Q�S0���T��   ��Gt61���[^_]Í�    ��    �B����   �83��   ��$��*	�v �P�S�x t��P�S�x�W���1w����$�h+	���&    1҉��W�������   P����M������[^_]Ív ��'    �P�S�x �Z����P�S�@��C<3�E������$�0,	��@���P�����t& �   닉���'    �C�R�����	����S�: ������z�{�:_������h��D$    ����'    ��������1�<$u�z  �v ��'    �7��t<$t��9�|������M���{)�����{������L$����  ���>   P����L���D$�����_���������=   ��j �L$�L�����@����t& �����������   j ���L����������&    ��'    ���Y����Ɖ�� R������   P���^L�����������    1҉�����������   j ���4L����������    ��    �x ��  �P�S�xn��  1҉����������H   j ����K�����n����v   ���vS�����X���1҉��u��������   j ���K�����6��������������   j ���K�������������������   j ���nK����������������ƍC�eP����������S�:_��������؉S�d����C0����V�   ���K���������h   ���R���������1҉����������   j ����J�����j���1҉��uR�����W���1҉��dR�����F���1҉��c��������   j ���J�����$������q��������   j ���~J�����������؉K0���������	   j ���VJ�����������
�؉K0�q��������
   j ���.J�����������O��������   j ���J�����������-��������   j ����I�����n��������������   j ����I�����L����G<St|<_tq<$�6����$   �S;S}j�C�4R���S����tW�H�{��� ?   ���{�r���f��D$����1҉����������G   j ���KI����������.   땹/   뎃C������    ��    UWVS���p���L��  ��T��  ��s���&  ��f��   �B�<	w6���������w  �S�ƀ:I��  ����[^_]�����������������o�W  ��t����  �~l��  �����������   � ��1��   ��2�\  ��3�  �C�8_��  ���0�����P��5   ���>H�������k����t& �~pu��F�C�~T�Z  ���N������  �S;S��  �K�4R���S�4�����  �   �F��������'    �F<r��  <p�+������؉s���������I   j ���G�����������f��E��7	��D$�@�֍H�K0�   ���������8��>  �D$�@����  ��  ���L  �E� �xc��  �؉T$�����T$�D$�(6	�   ����9  �7	�   ���t�7	�   �����  �������ƋC�8I��  ���7   ��V�L$�F����$�6   ���F������������1�����  ���E   �؉s�t��������0   P���rF�������������&    ��1�[��^_]Ít& �~n��������s�U����t& ��'    ��[^_]�����t& ��[^_]�DL���t& �E��������N  1҃��������u��.6	�   �����  �:n�q����B<at<w�a����_   ��襬���Ɖ�������S���<E�I  <p�q  <i�,����zl�"������[��������:   P���iE����$�9   ���XE����$�8   ���GE�������t�����    ��'    ���I�������   P���E�������D�����    ��'    ���؉s�#����Ɖ�������S�ǀ:I�Z  ��P��   ����D�������������1��s�����v ���H�������4   j ���D��������������E   �C���i����$����t& �<mt<p�
���:B�����C�8_�J  ���%��������7   P���3D���$������t& ��'    ���I�����P��������9����s���i�������������������������Ɖ�������ǉ������W���f��E   ��贪�����������    ��'    � �H���v��c<�j����؉T$�����T$�D$�e�����蛌�������   P���iC���$�������:�����������1��S��������_�������   P���-C�������S����zi��������؉S�E   ������������C������i�S����X�������'    U��WVS�Á�  ��d������`�����_��  �   �޿�4	�����1�8�u-�C<_��\�����<.��������M  ��\���$�@  ����\���S��  �����������l���ǅt���   ��p���� ����x���ǅ����    �����������   ���ǅ����    ǅ����    ǅ����    ���ǅ����    ǅ����    )�ǅ����    ��\�����)ă���|�����������  ��  ����  �{_�S��x���u
�{Z��  ����l���R��\�����  ��\�����������A��1҃�������j ��B�NA����x����Ɖ$��  ؃���x���� ���?  ���7  ��d����Uԉ��E�    �E� ���E�    �E�    �������E���`����E�    �E�    �E�    �E�    �E��E��E�    �E�    �E�    �E�    �E�    ��D���EԋM��E�    �ȍ�   ���)č�   �M�������U̺   )ĉ؉e��K���E�����Ƅ���� �u�PS�U��U���1������e�[^_]��C	<I��t
1�<D�����1��{
_������������������xZ�   �9����{�����_t%�e�1�[^_]Í�l��������Ƌ�x���� �����{ZuՍ�l������   ��x������S�����t�����u��x���� �Z�����x����<.�I����B�H�����   <_��   ��0<	w����<.u3��C��0<	w'�C�K�XЀ�	��wߍt& ����HЀ�	v�<.tΉى���x���)��?������K   P����>����x����ƃ��<.�l��������B�Z�H���w�����H���v�<_t��d�����l�����1҉�x������Q����5�����    ��    UWVS���D$0�t$4�\$<��t��t%�L$8��u����   �����1���[^_]Ð�t& �� 3�$    �D$    �D$    �D$    �E�������   �T$�<$�   ��Dl$��tV����   ��W�9�  ���T$8;sZ����PWV�V�  �<$���;�  ����tk�    ����[^_]Ít& ��'    ��t��tw�����1���[^_]Í�&    ��V���  �D$H���(뭍�    ��    �D$8��t��D$8�(둉����������'    ���t$譎  ����u�1�뚉���'    �����1�������v ���D$�T$��t!��t�L$�$�����������Ð��&    �������f�f�f�f��UWV���T$,�|$ �t$$�L$(�҉|$�4$��u=9���   �ɉ�u�   1���ŉ�1����Ɖ������^_]���������������;$w{�����   �    �׉�)�������	��<$���T$��D$�D$����������	ǉ��t$�Չ��d$9Չ$r�T$����9�sf;,$ua�G�1����^_]Ív 1�1����^_]Ív ��1�������^_]���������������;L$v1�;$�'����   ������t& ��1�����f�f�f��UWV�� �D$4�L$0�|$8�ƉD$�D$<�L$�|$�L$�t$����u9�vZ�ȉ�����1҃� ^_]É���'    9�w\���ud�l$9l$��   ;D$��   �D$�T$�� ^_]Í�    ��'    ����u�   1����ŋD$1�������덐�ȉ�� ^_]Ð�t& �    ��)���ǉD$�D$������D$	щ��L$�������D$�����ǋD$��щ����	��t$�t$����d$9щt$�׉�r
9D$s9�u�׉�+t$|$�ʉ�D$)�����L$�����	���� ^_]Ð�t$)�ƉL$�t$�����f�f�f�f�f��UW��V1�1ɍ�&    ���P��փ����	���x��w��@t	�������	׉} ^_]���������������U��WVS���O(  ��T ��<�}9։U�Ǉ�       ��   �E���   �}�@`�E���GL9���   �E��E�    �UЉEĉ���x�}ԉփ�����@t+����tt������   ��/�	  ����������t& �M��?���   �U�����   ;E�s'�}���   ���}Ћ}�O`�ʉM���WL9��x����e�[^_]É֋U�1���?1ɉ����Eȉ��EЍ�&    ���r���������	ǉ���x��uЋM�����   ����x����u�Mȍ��B   �:�a�����t& ��?����w�}�D�    �E��>���f��E��4�������  ����  �^�  �u�1�1ɉ׉���'    ���V��Ѓ�����	Ǆ�x���u�~h������}���   �����t���p�� �M���  v��MЀ�@��  ��P�$  ��0u��u�vX�uȉ���P�n  �������f����ҋ��P������}�P�����   UЉ��   �[����}�P�����   UЉ��   �<����}�����   �P�UЉ��   �����U�1�1ɍt& ��'    ���z���������	Ɖ���x��1҉u�1ɉƉ׍v ��'    ���V��Ѓ�����	Ǆ�x�����}�u����   ����������A   ������u�1�1ɉא�t& ���V��Ѓ�����	Ǆ�x�����j����M�D�    �Z����u�1�1ɉא�t& ���V��Ѓ�����	Ǆ�x�����*����M�D�   �����u�1�1ɉא�t& ���V��Ѓ�����	Ǆ�x����������u�D�    ������u�1�1ɉא�t& ���V��Ѓ�����	Ǆ�x��1�1��}ԉ�&    ��'    ���z���������	Ɖ���x�ЋUԃ��u����M���B   �2�a����}������a  ���   �}��ǹ)   �u�}���   �E��.����E�)   �}���   ���}��E����   �E������U�1�1�f����z���������	Ɖ���x�E��1�1ɉ��   ���׍t& ���V��Ѓ�����	Ǆ�x���}�����   Ǉ�      �����u�1�1ɉ׍t& ���V��Ѓ�����	Ǆ�x���u���   ǆ�      �[����u�1�1ɉ׍�    ���V��Ѓ�����	Ǆ�x���u���   �%����}�E�1�1ɉ��   Ǉ�      ��    ��'    ���z���������	Ɖ���x���������U�1�1ɍ�&    ���z���������	Ɖ���x���U�w�E���@   ��U�1�1ɉ���'    ���z���������	Ɖ���x����j����U�1�1ɍ�&    ���z���������	Ɖ���x�ЋU��-����}���   �U���#������A   ������U�1�1������������������z���������	Ɖ���x�}�ЋUĉ��   ������u�U����   ǆ�      ���   �����UċE������u�U����   ���   �����U�1�1ɐ��&    ���z���������	Ɖ���x��1҉u�1ɉƉ׍v ��'    ���V��Ѓ�����	Ǆ�x�����}�u����   ���������A   ��
����U�1�1ɍ�&    ���z���������	Ɖ���x�ЋU�������}���   �U����������A   ������U�1�1������������������z���������	Ɖ���x���U�w�E���@   ��U�1�1ɉ���'    ���z���������	Ɖ���x����:����E�1�1ɍ�&    ���p�������	׉��x�}�1�1����p�������	׉��x�u���   �uԃ�������M�ߍ��B   �:������P��1Ʌ�t�}��uȉ�Du�����   �ыu���   �����P��	���E�    ������P��붋Eԉ�1�1��M��׉���P��փ����	���x���}�뇋UċE��1����U��t����P���h����Uԃ�����B�
�t����u�v\�u��f����u�vT�u��X����
�Q������   �D$���������t& UW�z��VS�����1�)���L�    ���   ǂ�       ����G  ��J �Fh    �FP    �FL���l  �~`�ՍVT�t$��R�����|$�D�P��2  �D$$�������8  �F\�����   �ȃ�+A�D$�ǃ�	�D$P����  ���	e�D��  �L$�y�p  1�1ɍ�    ��    ���x��������	։���x�T$8���   1�������ƋD$81ɉ��   �D$�x��   �v ��'    ���V��Ѓ�����	Ǆ�x鉽�   �D$ƅ�   ��D$    � <z�e  �|$�L$<�L$ ���!�t& <Rtl<Ptx<S��  ƅ�   �������   <Lu�������   ������'    �   ��L[^_]Ív ������   �l�����������������������   �f��<��D$tu��p< �D$�  ��  �D$<@�  <P��  <0uG�D$�@X�D$(�|$P�F�D$$��  �D$��<w���������������.  <�&  藻  �t& ��'    �D$����  ���L$�U�t$�T�m������   ��<���  ��<��  ��  <��  <�   u�t$���    ��  1�1ɍt& ���V��Ѓ�����	Ǆ�x����   �<��D$��  �D$��p< �D$�F  �*����D$<@�C  <P�K  <0�����D$�@X�D$�|$P��  �D$��<���������������������'    �|$�
h����������|$���   ������t& ��'    1�1ɍ�    ��    ���V��Ѓ�����	Ǆ�x�>�|$ƅ�   �D$����|$�S������&    �D$���p����   �����v ��'    �V��1���t$�|$�D$(DD$$Ѐ|$ y� �t& ��'    ���   �����V��	�Ä�������   �R����V��먋t$$1҉|$,1ɉ׍t& ���V��Ѓ�����	Ǆ�x���|$,�t����T$ �D$$������T$<���\����V���P�����V��1���t�|$Et$��Ȁ|$ y� ��    �L$�։AP��D����L$�U�t$�T���������1��t�����V���1��|$ ��1ɉt$�Ǎ�    ���r���������	ǉ���x���t$�|$ �e�����V���X����T$<��� ����D$<���@�����V���3�����    ���   1�<��D$�G������B����t& ��t<������D$(    �;�����&    �F����p� �P����D$�@T�D$(�����D$�@\�D$(�����8������x ��������u����   �����   �x���������������V������D$�@T�D$������D$�@\�D$������D$    ������    ��'    UW��VS�  ��qC ��<  9Ջ�$T  �T$�D$0sx�D$(�D$   �D$��t& �0�x�N�������   �ɋ��������፴&    ��'    �l$�p����    ��?w{�}�t�0�|$;D$r��D$��tb�D�,��<  [^_]Ív �p�l$��	�čt& �F���8��$P  ��3�  ��$P  �Ac@�4�t�|l ��  ����  ��t& �W�  �t& ��'    ���y�������'    �p�l$���P����p�l$���@����p�l$���0����p�l$��� ����t$��t��������t�0�t$��  �L  ��#�  �����  �� �a����t$����������t& �x������A�����p�� �T$�U  �!  �T$��@�g  ��P�  ��0������$P  �vX�t$�p����P�t$��  ������������ҋ��������⍴&    ��'    1�1ɍ�    ��    ���W��Ѓ�����	ń�x���������$P  ��$P  ��+�  �Bc@�4�t�|*l u���a����6�l$��������t& �T$���U����V����9�����$P  ��3p  �Gc@�4�t�|l u�������6t$(�e  ��    �D$��������P����t�0�L�0�t�0�L�0���f�����    �l$�H�P����L$(9������)ȋt�0���'�����&    �P�D�#����v �t$����������P���L�0�t$��������������v �D$���S����h����L�,���t�0�<����ҋ�����������&    ��'    �D$�������H��P����t�0�l�0�t$�t�0�t�0�t$�t�0�l�0���s����v ��0�l$���R���f��D$��������t�,�ŉ��7�����&    �T$,�������t$,�l$�������&    ��1�1ɍv ��'    ���x��������	։���x��Đ�t& 1�1ɍ�    ��    ���W��Ѓ�����	Ƅ�x�T$���>������%�����$P  ��3�  �Gc@��t�|7l u����������t$(�O����D$��������t�(�ŉ��V�����    �D$����������D$���F�����$P  �v\�t$�����p�����l$�����|$�T$DT$։���������6�������1�1ɍv ��'    ���x��������	։���x�t$�����p��
뙍�    ��tb���"����T$��������1�Ɖ�������t	��������D$    ��������l$����0���\�����$P  �vT�t$������D$�0���<����P�@<�q  �U  <t<������D$�0�������t$����������������	Ή������Ή�������������������������������1Ή������1�9����Ɖ�����!Ή����������Ɖ�����)Ή�������1����������1�9����Ɖ��r���1�9����Ɖ��b���1�9����Ɖ��R���1�9����Ɖ��B���1�9����Ɖ��2����D$�T$,�����t$,������p��������p��������D$1�1ɍ�    ��    ���h�������	։��x�����<�J����D$�0�������D$�0��������&    ��'    UW�    VS����  �Ì; ��   �|$0�D$�T$�|$���$�   @��   ��$�    ��   �D$�@c@t�@p �D$�@    �D$���   ����  ����   �D$1�1ɋ��   �v ���p�������	׉��x���8j �t$$�f����D$$���D$�t$�D$    �pH�t$��l�D$��~wl�F���0��������    ��    �D$@���>������  �D$�@H�b  �W�  �t& ��'    �D$�|$���  w܋L$��L$���D$���D$�D$���t����D$���    �D$��  �``����ļ   [^_]Í�    ��'    �1�1ɍv ��'    ���x��������	Չ���x���(�t$�t$$�D������|$�Gc@t�L$� �L$�|$���R����1�1ɍv ��'    ���x��������	Չ���x���(�t$�t$$��������L$���  ������|$��|$���������    ��    ����    uT�L$�D�0�Ac@�b����V�����    ��'    �|$�D$�Gc@t�L$� �|$�L$����������'    ���G�����$�   @���  �D�0�C������$���� �3�����    ��'    �D$���   ���������$�   @���  �T�0t'���    t�D$��   �T$�k����v ��'    ���������֍v �H`   ��ļ   [^_]���$�   @�D$,tƄ$�    �D$,�D$@�����t& ��'    UW�x��VS����Ɖ�)����   �     ���@|    1����|$�F`   @��  �í7 ��$�   ���FL���X�����u���   t���  �~   �U�  ����'    ƃ�  ƃ�  ƃ�  ƃ�  ƃ�  ƃ�  ƃ�  ƃ�  ƃ�  ƃ�  ƃ�  ƃ�  ƃ�  ƃ�  ƃ�  ƃ�  �Fc@�l$t�Fp �D$��Ǆ$�      Ǆ$�      Ǆ$�       �F���!�����$�   �FL���   [^_]Í�    ��    WV��S����
  �Ð6 ��������   �|�t<���Fc@���  ��u��t1�8�  ��    ��    �|l t�[�VL^_�f�[�FL    ^_Ð�t& ��㍶    ��    UW��VS���O
  ��6 ���   �l$�B���$�   ��t)����VW���w�7�T$$Qj�Ѓ� ��tU���T$u1��uX�����������v����V`�NH��)�9O��������t����   �   [^_]Ít& ��'    ���   �   [^_]��G�  �t& ��'    UW��V�Ɓ��   �@�l$�D$�F�D$�c�����������������t$WV�v�6j
j�D$$�Ѓ� ���}   ��$�   ��t��WV�v�6j
j�Ѓ� ��tj��uU����<������������t��u:��u��D$���t$WV�v�6jj�D$$�Ѓ� ���T$u�Ё��   ^_]�f����   �   ^_]Ð���ލv ��'    UW��VS�  ��a4 ��,�Bc@tV�zp tP1��T$�v ��'    �|l �|� �L$�|$�4�u ���|l ��tL��tH���  ��   ��  ��t& �r��u����  �BHu��Bc@�D$t�Bp �D$�B농�    �����D$�T$��t.9t$t(���  ��s[��t��T$��   �
��   f������D���1��Ec@�T$uh�M��to��,[^_]É���'    �T$�2�Ȑ��&    ��T$�
�L7��L��T$�J�T$����L$)ʉ�)���|$���닍t& ��'    �}p t���,[^_]��Bc@���  �Bt�zp u�������� +EHBh��,[^_]��t7��T$f�t��0���VS��  �õ2 ���T$�L$���Ac@���  ��u��t�d�  ���&    �|l t��[^Ív � ��[^Ð��&    �D$�@HÐ��&    S�  ��F2 ���D$�T$���Bc@���  u����t.���  ����'    �|l t�L$����[Í�    ��'    �L$���[Ð�t& �D$�@LÐ��&    �T$�L$�B`����BLÍ�    ��    �T$�D$�PLÍt& �D$�@PÐ��&    �D$�@\Ð��&    S�  ��v1 �� �D$P�D$,��P�  ����t�D$��[���������������1��荶    ��    �D$�@XÐ��&    �D$�@TÐ��&    UW1�V�    ��@  �狴$T  󫋄$P  ��$�   �D$`   @�����D$L����������   ��$   ty1������'    <t�D�    ����t�D�<�D\u��ωD�����u勄$  �F��$  f�FX��$4  f�FZ�D$h�F��$<  �F��@  ��^_]Á�@  1�^_]Ð��&    ���������������U��WVSR��(���P�������U�����  �u�� ���������$����    ��󥍵(����J�t& ��'    ��ul�EЅ�t'�}����$����u�w�7jj�Ѓ� ��tS��u>��$������������$������D�����u��   �]�u��}������������������   �]�u��}��ËE��������$�����$����� ����@    �������)��ȋM�A�E�    ��������u���$����� �����������������W������������|5���L�E�U��]�u��}��m ��Í�    ��'    U��WVSR������P�U��h�������   �u�����������U�E�    󥍽h������B�E�щB�����������t�]�u��}��Ë�������������}���PPW�u��������|5���L�E�U��]�u��}��m ��Ív ��'    U��WVSR������P�U��h����   ���- ��   �u��������������E�������    ���������H��u������t�u�  �E�1����싕���������������}���PPW�u��>�����|5���L�E�U��]�u��}��m ��Í�    ��    U��WVSRP�o  ��/- ��  �E�@��tM���������U�u��h����������������    �E��󥍽h�����������t,賠  ��&    ���u�������]�u��}��Í�&    ���������3����}�����W�u��b�����|5���L�E�U��]�u��}��m ��Ã��T$�B��t��Rj�Ѓ���Ív U��WV�������U��\  �u���B�����8������������$����uV�U����u*��t:���������]�������������������tɅ�tōe��   ^_]É���'    �e��   ^_]Ë$�UW��V1�1ɍ�&    ���P��փ����	���x��w��@t	�������	׉} ^_]����������������L$�T$�B9A�R�9Q�   G�ÐUWV���T$�T$$�$�|;|$(|D�   �D$ ���,��D$ ���u �<��7�t$�D$�Ѓ���yg�U ���|69|$(�E ~S��w9t$(~��D$ ��    �T$���L$�l��D$$�4��u �t$�D$�Ѓ����L$�T$x��뀍�&    ��^_]É���'    L$ ���^�����t& UWV���D$�D$ �T$�p�h��������t*��    ��    ��VW��U�T$�D$����������u���|$ ��~1��&    �T� �G���W�D� Vj U�T$�D$��������uփ�^_]���������������S�������) ��<�t]����tCv!��t ���   u"��[Í�    ��'    ��u���   [�f��g�  �t& ��'    ���   [Í�    ��1�[É���'    S������V) ��<�t=��p< tFv<0u �B��[Ð��&    ��t<t���  �v <Pu�    ��    ��1�[É���'    �B��[Ð��&    UW��VS�!������( ��,<P�T$��   ����<��   �����H��������t& �D$@��p��t����p<�D$DD$@���y��D$D���,��[^_]É���'    �D$@��p뾐�t& �D$@��p뭍t& �D$@�T$�����T$��딍t& ��'    �t$@1�1ɉՍ�    ���V��Ѓ�����	ń�x���[���f��D$@��p�J�����Ǜ  �t& ��'    �D$@�p�D$D���������,��[^_]ÐUWV���l$ �E��f�������B������ǍD$��P�D$0��P������XZ�E�T$f��R�L$4���QR���v����D$9D$�   �t$�9t$G� ^_]Ð�t& WV�x	S���o�����/' ��W��  ���~�L��   �~	zt1���[^_Ít& ���y� x��T$���,����~����   ���z� x��~
�t& ���z� x��F
�t$<Ru�I����'    <Lu������<Rt/<Pu���J��V1҃�Q�����������<Ru؍�&    ���[^_Í�    �9��   �G����y �=������-������a������&    UWV�փ�0����J  �ōD$,�D$    �D$    �D$    1ɉD$�v ��'    �F����   �~)�9���   ������=�   �D$��   �D$��D$�R����D$�E��f���f�����   f����9D$t�M�F���t$ P�T$$�D$�����D$�������������w��    �   ����D$,����t�D$;E s�E ����t����/����D$��0^_]Ít& �T$f%���	�f�E�r�������'    �D$�D$�[���f���0�����^_]��D$    뫍v ��'    UW��V��0�@�t$@�T$��f�������<�����D$�D$,�D$    �D$��u@��   ��    ��'    �V��t�D$� ��t�P�J�H�t���t�����   �V��t��Et&�N)�9L$t�ȉL$���������������D$��t������ȍF�t$$P�T$ �ȉL$(������L$(���������������w��    �   ����T$,�P�����t����g�������'    ��0^_]É���'    UWV�։� �$�@f�D$f�����������.�D$�D$�D$    �D$��uB��   ��    ��'    �F�V���D$�T$t�L$0)�9���   ��t�����   �V��t�$�@t'�n)�9l$t�������$���������l$�D$��t�������F�t$P�T$�������ZY�����T$$RP1҉��������������������w��    �   ����D$���S����L$0�T$)�9��A����� ��^_]Ð��&    �� 1�^_]Í�&    UWV���|$$�t$(�G+G��������T$ ����������T$RW�������F+F�������T$0��������ZY�T$RV��������D$9D$�   �L$�9L$G� ^_]Í�    UW��VS������á! ��L�@�T$���   ���  �uf����1  �u1�F���D$�D$9�vV�L ��D��p9t$�P�T$��  �|$�.�t& ��'    �)�D$��D��p9t$�x�|$��   ��9�r�1���L[^_]����������������M���ɉL$(��  ���  �u���tA�������'    ���ǅ���  ���z������u��  �E    f�E���  �E�D$9E �v����E��������  �u����U����|$�v ��'    ����W���������3��������u��#�����    ��    �|$t$9t$�����j�L$����f��E�D$$�@���D$������D$8�D$    �l$(�D$ �D$4�D$�/��    ��    D$8;D$�  �E�D$�L$9L$������l$l$�D$$��|��G+G�@����T$(�ȉƉȉL$���	����W���t$$R�L$(���a���ZY�t$(P1҉��Q����D$D��;D$�p����l$�|����U�����������D$(�k����L$(��%�� 9��]  �e�  �D$(���^����D$(���4�   V��O  �D$H�������9������@    V�O  �D$L����t�@    �E��  �u����<  �L$8�ύ�    ������P�����������u�D$8�D$,�|$,��t�D$,�L$(;H��  �E������uf�E���������D���DǋD$<���D$��  �L$,�A���D$ ��  �ȍ��  �|$���D$$    �D$�L$�ωƍ�    ��'    �D$$�L$�|���;D$ �D$$�?  ;t$�)  ���#��t& ��+D$D$�x;|$�@    �  ���7�vU�D$(�Ѓ���x̃�뗍�&    ���U���t$��������L[^_]ËEf����ǉD$�����D$������o�D$$��������1Ƀ��ΉD$(�D$8�D$ �D$4�D$�"����'    D$8;D$�;  �w9�������D$�<.����L��t$$�A�L$P�T$4�D$(����ZY�t$(P1ҋD$8�����D$D���L$;D$v���먍�&    �|$������1�1�1ҋ|$�t$�L$,�l$���    ��    �t�����;T$ t�t����t�u�l$�t��u�t$�ڋL$8�|$�l$�T$<�t$�L$�L$,�A�D$�p�D$�@B9D$(��  ����R���\����D$L�L$H�D$4�@�D$0������   �Q���|$�l$�͉D$�א��&    �l$ �T$$���D$ �D��D$��   �������t& ��'    �D��T$�����D�t~�u����t$�t��t$$�D$,�Ѓ���ω���ǋL$ �T$�l$����ɉT�u��D$$��l$�@A�D$<�D$$���t$0�R  ���D$8�U��E�M�X����t& ��1�롉|$(��������D$D�u��������D$H�D$<���O����������������U�������  	ЉE�����ʋL$�a����������t$8��������l����D$,�T$1��D$1��E����|$,�������  f�S�T$�r�����2 �D$��t<�
��t6�L$�P��  �@    � �����H�L$f�P��  ��  �H�P[Ív ��'    �T$�D$�#  ��� ��t�: u��f��P��  �@    f�P��  � �����@    �@    ��  �PÉ���'    VS������u ���t$���tC��j�WJ  ��  �@    � ����f�P��  ���@    �@    �p��  �P��[^Í�    ��'    �D$�T$�S  ��� �P�T$�@    �@� �����P�T$f�H��P��  ��  �PÐ�t& �D$�T$�  ��� �@    �@f�H��P��  � �����@    �@    ��  �PÐ�t& S������f ��j�UI  �T$ �@    �@f�H�� �����@    �P��  �@    ��  �P��[Ív ��'    VS�E����� ���L$ ����   �����   ��  ��t9Ju�   ��    9HtK�B��u�   ��tH��   ��p9tY�P�@��t/�@u�9Hu�H�
��[^É���'    ����t& ��'    �G�  �t& ��'    ��1�[^Ð��&    �H���
�p�D$�UN  ���D$��[^ÉЍ�  두�t& �����t& ��'    S�F����� ���D$���t��P������$��M  ����[Í�&    ��'    UWVS������� ����   �|$0��u�   �t& ��'    �v����   9>w�������������t{�F�|$4��F�G�Ff���F��t�E+E�����������������T$R�UR���F����D$�|$D���G����[^_]Í�   ���&    ���M�*uN��  ��tՋE����  ���;�����   ��tËu ;1v뺐��&    ;1w��Q�I��u���M�*t�����.����$�U����E�E��E���Ph  �  ���E���U���j jj �u�2  ����U���j j�u�u�  ����U����E�E��E���Ph  �  ���E���U����E��Ph  �  ���E���U�����h   �u�   ����U����E�E�E�E��E��Ph  �Z  ���E���U����E�E�E��Ph  �5  ����U�����j j j �u�u�f   �� ��U�����j �uj �u�u�F   �� ��U�����j j �u�u�u�&   �� ��U�����j �u�u�u�u�   �� ��U���(�E�E��E�E�E�E�E�E�E�E��E���Ph  �{  ���E���U���(�E�E��E�E�E�E︐0�E�E��Ph  �A  ���E���U����    U�����j h  �  ����U�����j j �u�u�u�G   �� ��U������uj �u�u�u�&   �� ��U�����j �u�u�u�u�   �� ��U���(�E�E�E�E�E�E��E�E�E�E��E���Ph  �|   ���E���U�����j �u�   ����U����E�E�E�E��E��Ph  �9   ���E���U����E�E�E�E��E�E�E��Ph  �   ���E���U��S�E�U��̀[]�U����E�E�E��Ph  ��������E���U���(�U�E�U�E��E�E�E�E��E�������E����	ЈE��E������ �E����	ЈE��E�����E��E��Ph	  �_������E�������U������u�#   ����u�E��0��	w�   ��    ����U������u�j   ����u���u�  ����t�   ��    ����U��} x�}�   ��    ��]�U��} ~�}~�   ��    ��]�U��}`~�}z�   ��    ��]�U��}~�}~�   ��    ��]�U������u��������t���u���������u�   ��    ����U��} t�}t�}
t�}t�}	t�}u�   ��    ��]�U��}@~�}Z�   ��    ��]�U��}/~�}9~�}`~�}f~�}@~�}F�   ��    ��]�U��}@~�}Z�E�� ��E]�U��}`~�}z�E�� ��E]�U��]�U��    ]�U����x   �L���E��������E�P�E�P�A�  ��������t5�E� ��P�@�  ����P�������U�E���RP�eN�����E����h�W	���������u��5�  U�����h�W	j �^�������j j��l  ���G~  ��U����  ��U����E�    ��E��E��?������t�l  �E� ��u�U�   ���t�   ��    ��u��    ��U����E�  �E��E�� ;Ew�E���E��@�;Ev�E���E��@�E��}� ����t�    �����U����E�  �E��E� ;E�w�E��E�@�;E�v�   ��E��@�E��}� ����t�    �����U����   ��[��t��h�[���������[����   �E�   �E�E�   ��v9�   �   ��!Ѕ�u&�   ����u�E���#E���u�E��#E��t�e�  �E�[�E���[��[������[    ��[   ��[�|]��]    ��j �߈  ��5UUUU�E�M��e����[�E��    ��[�   ��U�����[��u	�������t��}�t�E�������E�E���t���t���t>�K�E���[�   �A��[;E�w�E��#E��u�E���[�   ��    ��E���[�   ��    ��U��WS�� �E�ø    �
   �߉�󫡄[��u	�B�����t��E���  ����t,�E���  �   ���t�E�  ��P��������u�   ��    ����  �E�@����  �E�   �E�@�   �   ��!ʅ�t"�   �   �   ��!�)Ѻ   ��!���    �   �   ٍY��   ��!�Ѻ   ���Z��   ��!��ЉE��E��E�E�  �E���   �E��E� �   ȉ��   ��!ȅ�t+�   �E� �   ؉ø   ��!�)��   ��!���    ЉE��6�E�@����E��E�E�E�@����u
�E�E��E��E�@���E�E� ;E�w,�E��E�@�;E�v�E�@;E�t�E�@�   9�u��E�@�E�}� �)����E�U��E�U�P�E���  +E�E�P�E���  �E�P�E���  +E��E�P�E�U��P �E�P�E�P$�E���  ����t�E�  �    ���E�e�[_]� U��S��$��[��u	�������t��E���  ����t,�E���  �   ���t�E�  ��P��������u�   ��    ����  �E�    �E�    �E�    �E�@���i  �E�  �E�E���  �E�E���  �E��E�@�   �   ��!ʅ�t"�   �   �   ��!�)Ѻ   ��!���    �   �   ٍY��   ��!�Ѻ   ���Z��   ��!��E�)ЉE��   �E��E� �   ȉ��   ��!ȅ�t+�   �E� �   ؉ø   ��!�)��   ��!���    ЉE��&�E�@����u�E�@���)E�E�@���E�E� ;E�w,�E��E�@�;E�v�E�@;E�t�E�@�   9�u��E�@�E�}� �9����E���  ����t�E�  �    ���D���u�h`Y	P�k  ����D���u�hzY	P��j  ����D���u�h�Y	P��j  ���]���U��� �   �   Eк   ¡�[ЍP���[��!ЉE��E���  ��t7�E���  �E�ЉE��E���  ;E�s�E���  ;E�s
�    �)  �E�;E�  �E������}���  �   �E�Љ¸   ��!Ѕ�t)�   �   �E�ȉ��   ��!�)¸   ��!���    �E��E�+E�   )ЉE�U�E�ЉE�E�U���E�U�P�U�E�к   �P�E�P�E���@    �E�@��t�E�@;E�v	�E�U�P�E���  �E�E���  �E���  �E���  9�����t�E���  �E���  �   �E����    ��U��� �E�@����E��E����w
�    �)  �E��;E�w�E�+E��[�9�w�E�  �E� �E��U��E�к   ЉE��   �   Eк   ¡�[ЍP���[��!ЉE��E������}����   �U�E�ЉE�E�+E��   )ЉE�E�U�P�U�E�к   �P�E�P�E���@    �E�@;E�v	�E�U�P�E���  �E�+E�E���  �E���  �E���  9�����t�E���  �E���  �E���    ��U��S���   �EЉ¸   ��!Ѕ�t)�   �   �Eȉ��   ��!�)¸   ��!���    �E��E�E�E�)E�E�U�P�E�U�P�E���E�P�U�Eй   �   ��!ʅ�t"�   �   �   ��!�)Ѻ   ��!���    �   �   ٍY��   ��!�Ѻ   ���Z��   ��!�ʉP��[�E�P��[]�U����E�    �3�E������    �EЃ��E��E��U��P�E��P�E��P�E��}�v���U��S��   �   �EЉ¸   ��!Ѕ�t)�   �   �Eȉ��   ��!�)¸   ��!���    �EЉEк   �EЉ¸   ��!Ѕ�t)�   �   �Eȉ��   ��!�)¸   ��!���    �EЉE�U�E�)ЉE̋UЋEЉEȋE�+E�E��E���EЉP�E�@;E�u6�E�P�E�E�P�E�@�EċE�UȉP�Eă��EȉP�  �E�@;E�uC�E�P�E�E�P�E�@�E��E�UȉP�E����EȉP�UȋE�E����  �E�@������  �E�@����E��E�������   �E�@�E��E�@�E��E����E��E������    �EЃ�;E�t�E�@;E�w�E��@;E�u�   ��    ������   �E�;E�u�E��E��   �������!E��c�E������    �EЃ�;E�t�E�@;E�w�E��@;E�u�   ��    ����t�E��U��P�E��U��P�
�t  �t  �p  �E�E��E��@�E��E��@;E�tb�E��@�E��E��@�E�E�@;E�w�E��@;E�u�E�@;E�u�   ��    ����t�E��U�P�E�U��P�   �-t  �E����E�E� �E�}� u�E����E�E� �E�}� t�   ��    ��tg��E�E�E� �E�E���E�E� ��u�E���E�E� ��t�   ��    ��u��E�@;E�������t�E��     ��s  �}� �E  �E��@��L��    �EЉE��E�� ;E�u9�E��U��E�� ������t\�E�P�E��@�   �������!E�P�9�E�@;E�������t!�E��@;E�u�E��U�P��E��U�P���r  �}� ��   �E�@;E���������   �E�U��P�E��@�E��}� ����t,�E�@;E�������t�E�U��P�E��U�P��r  �E��@�E��}� ����t,�E�@;E�������t�E�U��P�E��U�P��@r  ��9r  �E�E�E�E��E�@����E�P�E����EȉP�UȋE�E���E�������   �E����E��E������    �EЃ��E��E��E��E��E�����Ѓ���u�E��E��   �����	E��(�E��P�E�@9�������t�E��@�E���pq  �E��UȉP�E��UȉP�EȋU��P�EȋU��P�E  �EȉE��E����E��}� u	�E�    �C�}���  v	�E�   �1�    �E���)Ѓ��E��E�� �E������E����ЉE܋E܃�L��    �EЉE��E��U܉P�E��@    �E��P�E��P�E�P�E܉���Ѓ���uG�E�P�Eܻ   �����	E�P�E��U���E��U��P�E��U��P�E��P�E��P�S  �E�� �E؃}�t�    �E���)Ѓ�����    �E������EԋE؋@���;E���   �    ���Eԉ��������    �E�Љ�|����eԋ�|���� ��t��|���� �E���   �E�@;�|���������t.��|����U���E��U؉P�E��U��P�E��P�E��P�   �o  �E؋@��x����E�@;E�w�E�@;�x���w�   ��    ����t<��x����U��P��x����P�E؉P�E���x����P�E��U؉P�E��@    �
�o  ������   �E�ЁĄ   []�U��S��   �E�@�E��u��u�A������E؋E؋�E؋@ЉEԺ   �   ЍP��   ��!ЉEк   �E�к   к   )E�ЉE̺   �E�Љ¸   ��!Ѕ�t)�   �   �E�ȉ��   ��!�)¸   ��!���    �EȋŰE�ЉEĸ   ���P��   ��!E��;E�v�E���EĉE��E��E��   �E�ЉE��U��E�ЉE��E��E��E�    �   �   ��!Ѕ�t"�   �   �   ��!�)¸   ��!���    �   �   ʍJ��   ��!�¸   ���H��   ��!�E)�P�u�u��������EЃ��E��P�E��U���  ����  �H���  �H���  �P�E�U���  �E�U���  �E�U���  �E�U����  �E���E��   �E�P�E��E���;E�s�E��E����E�;E��(  ��ċE܉E��U��E�)ЉE��U��E�ЉE��E��@����E��P�E����E��P�U��E�E���E�������   �E����E��E������    �EЃ��E��E��E�E��E�����Ѓ���u�E��E��   �����	E��(�E��P�E�@9�������t�E��@�E����k  �E��U��P�E�U��P�E��U�P�E��U��P�   �E��E��E����E��}� u	�E�    �C�}���  v	�E�   �1�    �E���)Ѓ��E��E�� �E������E����ЉE�E��L��    �EЉE��E��U�P�E��@    �E��P�E��P�E�P�E����Ѓ���uG�E�P�E�   �����	E�P�E��U���E��U��P�E��U��P�E��P�E��P�.  �E�� �E�}�t�    �E���)Ѓ�����    �E������E��E�@���;E�t�    ���E����������    �E�ЉE��e��E�� ��t�E�� �E��   �E�@;E�������t(�E��U���E��U�P�E��U��P�E��P�E��P�t� j  �E�@�E��E�@;E�w�E�@;E�w�   ��    ����t3�E��U��P�E��P�E�P�E��U��P�E��U�P�E��@    �
�i  �����]���U��S��d�E������E�    �E�    ��[��u	�v�����t� �   �   ��!Ѕ�t"�   �   �   ��!�)¸   ��!���    �   �   ʍJ��   ��!�¸   ���H��   ��!�к   E¡�[ЍP���[��!ЉE܋E�;Ew
�    �	  �E���  ��t7�E���  �E�ЉE؋E���  ;E�s�E���  ;E�s
�    ��  �E���  ������  �E������E܉E�E�@��t�E�@��P�u��������    �EԸ   ��[��t��h�[�/������}� ��   ��j �qq  ���EЃ}����   ��[�P��E�!Ѕ�t!��[�E�ЍP���[��!E�)�E�E���  �E�ЉE̋E�;EvS�}����wJ�E���  ��t�E���  ;E�s/�E���  ;E�r!�E��P��p  ���E�E�;E�u�   ��    ��t�EЉE�E�E���   �E�@�U)¹   �   ��!ȅ�t"�   �   �   ��!�)��   ��!���    �   �   ٍY��   ��!���   ���X��   ��!�ȹ   �¡�[ЍP���[��!ЉE�}����w+�E��P� p  ���E�Eԋ�Eԋ@�9E�u�   ��    ��t�E�E�E�E��}����  �}���^  �}�����Q  �   �   ��!Ѕ�t"�   �   �   ��!�)¸   ��!���    �   �   ʍJ��   ��!�¸   ���H��   ��!�к   E�;E���   �   �   ��!Ѕ�t"�   �   �   ��!�)¸   ��!���    �   �   ʍJ��   ��!�¸   ���H��   ��!�к   E�+E�¡�[ЍP���[��!ЉEȁ}����w8�Eȃ�P�n  ���Eă}��t�E�E���E��؃�P�dn  ���E������}��t�E�E�E�E���E���  ���E���  �    ��[�}���  �}�����  �E������E������   ��[��t��h�[�������E܃�P��m  ���E���j ��m  ���E��    ��[�}����   �}����   �E�;E���   �U��E�)ЉE��   �   ��!Ѕ�t"�   �   �   ��!�)¸   ��!���    �   �   ʍJ��   ��!�¸   ���H��   ��!�E�;E�s�E��E�E��E��}����  �E���  �E�E���  �E���  �E���  9�����t�E���  �E���  �E�@����  �E�@��t�E�@;E�v	�E�U�P�E�U��  �E�U����  �E�U����  ��[�E�P$�E�@ �������u�[������}�[��   �   �   ��!Ѕ�t"�   �   �   ��!�)¸   ��!���    �   �   ʍJ��   ��!�¸   ���H��   ��!�E�)Ѓ�P�u��u��������	  �   �؉EЋ@����   )ЉEЉE��U�E�ЉE�)Љú   �   ��!Ѕ�t"�   �   �   ��!�)¸   ��!���    �   �   ʍJ��   ��!�¸   ���H��   ��!��)É؃�P�u��u�������L  �E�  �E��	�E�@�E�}� t�E��E�@�;E�u߃}� tp�E�@����uc�}� u]�E�P�E� 9�rN�E�P�E��E�@�9�s7�E�P�E�E�P�E�P�E�E�@��RP�u�g������   �E�@;E�v	�E�U�P�E�  �E��	�E�@�E�}� t�E� �M�U��9�u��}� tM�E�@����u@�}� u:�E� �E��E�U��E�P�E�E�P�u�u��u��u�"������   �u��u��u��u�J������E�@;Evb�E�@+E�E�P�E�@�E��E�@�E��U��EE�P�E�@�E��E����E��P�E���E��P�   �E���e�    ������2   �    �]���U��� �E�    �E�    �E�  �E��E��@�E��*�E�� �E�E��@�E�E��@�E�E��E��E��E�E��}� uЋE�@ �����E���U���(�E�    ��[��u	�<�����t��   ���P��   ��!�����;E��  �E�@����  �   �   ��!Ѕ�t"�   �   �   ��!�)¸   ��!���    �   �   ʍJ��   ��!�¸   ���H��   ��!��E�E�@;E�C  ��[�E�E�@+E�E�Ѓ��    �u���E�E��E�@��P�u�������E�E�@������   �}����v�   �+E�E�   ��[��t��h�[��������j �Xg  ���E�E��E�@�;E�u?�E��؃�P�2g  ���E���j �"g  ���E܃}��t�E�;E�s�U�E�)ЉE��    ��[�}� tI�E�@+E�E�P�E���  +E�E���  �E�@+E�E�@��RP�u�������}� u�E�P�E�@9�v
�E�@�����}� t�   ��    ��U��S��   �U�EЉE̋E�@�����*  �E� �EȋE�@����u�   �E��E�{  �E��؉EЉEċE�E�EĉE�E�@;E���������  �E�@;E�s  �E�������   �E�@�E��E�@�E��E����E��E������    �EЃ�;E�t�E�@;E�w�E��@;Eu�   ��    ������   �E�;E�u�E��E��   �������!E��c�E������    �EЃ�;E�t�E�@;E�w�E��@;Eu�   ��    ����t�E��U��P�E��U��P�
�{[  �v[  �p  �E�E��E��@�E��E��@;E�tb�E��@�E��E��@�E�E�@;E�w�E��@;E�u�E�@;E�u�   ��    ����t�E��U�P�E�U��P�   ��Z  �E����E��E�� �E�}� u�E����E��E�� �E�}� t�   ��    ��tg��E�E��E�� �E�E���E�E� ��u�E���E�E� ��t�   ��    ��u��E�@;E�������t�E��     ��PZ  �}� �E  �E��@��L��    �EЉE��E�� ;E�u9�E��U��E�� ������t\�E�P�E��@�   �������!E�P�9�E�@;E�������t!�E��@;E�u�E��U�P��E��U�P��Y  �}� ��   �E�@;E���������   �E�U��P�E��@�E��}� ����t,�E�@;E�������t�E�U��P�E��U�P��HY  �E��@�E��}� ����t,�E�@;E�������t�E�U��P�E��U�P��Y  ��Y  �H�E̋@����u:�E�U�P�E̋@����ẺP�E���E�P�U�EE��  ��X  �E�@;E��������\  �E̋@������  �E�@;E�uU�E�P�EE�P�E�@�E��E�U�P�E����E�P�E�@;Eu�E�@    �E�@    ��  �E�@;E�uC�E�P�EE�P�E�@�E��E�U�P�E����E�P�U�E�E���  �E̋@����E��E�E�E�������   �E̋@�E��E̋@�E��E����E��E������    �EЃ�;E�t�E�@;E�w�E��@;E�u�   ��    ������   �E�;E�u�E��E��   �������!E��c�E������    �EЃ�;E�t�E�@;E�w�E��@;E�u�   ��    ����t�E��U��P�E��U��P�
��V  ��V  �  �ẺE��E��@�E��E��@;E�tq�E��@��|����E��@�E�E�@;�|���w ��|����@;E�u�E�@;E�u�   ��    ����t��|����U�P�E苕|����P�   �<V  �E����E�E� �E�}� u�E����E�E� �E�}� t�   ��    ��tg��E��E�E� �E�E���E��E�� ��u�E���E��E�� ��t�   ��    ��u��E�@;E�������t�E��     ��U  �}� �o  �E��@��L��    �EЉ�x�����x���� ;E�u?��x����U���x���� ������t\�E�P�E��@�   �������!E�P�9�E�@;E�������t!�E��@;E�u�E��U�P��E��U�P���T  �}� ��   �E�@;E���������   �E�U��P�E��@��t�����t��� ����t5�E�@;�t���������t�E苕t����P��t����U�P��tT  �E��@��p�����p��� ����t5�E�@;�p���������t�E苕p����P��p����U�P��%T  ��T  �E���E�P�U�EE��E�@;Eu�E�U�P�  �,�E̋@����ẺP�E���E�P�U�EE��E������   �E����l�����l��������    �EЃ���h�����h����E܋E���l�������Ѓ���u�E���l����   �����	E��.��h����P�E�@9�������t��h����@�E���S  ��h����U�P�E܋U�P�E�U܉P�E��h����P�  �E��d����E����`�����`��� u	�E�    �R��`�����  v	�E�   �=�    ��`�����)Ѓ���\�����\���� ��\��������E���ЉE؋E؃�L��    �EЉ�X�����d����U؉P��d����@    ��d����P��d����P�E�P�E؉���Ѓ���u_�E�P�Eػ   �����	E�P��X�����d������d�����X����P��d�����d����P��d����P��d����P�t  ��X���� �Eԃ}�t�    �E���)Ѓ�����    �E�����EЋEԋ@���;E��   �    ���EЉ��������    �E�Љ�T����eЋ�T���� ��t��T���� �E���   �E�@;�T���������t@��T�����d������d����UԉP��d�����d����P��d����P��d����P�   ��P  �Eԋ@��P����E�@;E�w�E�@;�P���w�   ��    ����tH��P�����d����P��P����P�EԉP��d�����P����P��d����UԉP��d����@    �
�DP  �������8P  �Ĵ   []�U��S��   �E�    �E�؉E��E���E��}� u	�E�    �C�}���  v	�E�   �1�    �E���)Ѓ��E��E�� �E������E���ЉE�E�U��L���E�}� ������   �}�t�    �E���)Ѓ�����    �E�����E��E�    �E�@���+E�E��E�;E�s�E�E�E��E��}� ����t�U�E�@�E��    ���E������E�����E�}� t�E�;E�t�E��E��}� u�E��E���e��{����}� ud�}� u^�E�   ����Ѝ �E�   ��������	E�@!ЉE��}� t(�E���#E��E���E��E��E��E��E�U���L���E��>�E�@���+E�E��E�;E�s�E��E��E�E�E�@��t�E�@��E�@�E�}� u��}� ��  �E�@+E;E���  �E�@;E��������q  �U�EЉE��E�;E��������R  �E�@�E��E�@;E�tb�E�@�E��E�@�E܋E�@;E�w�E��@;E�u�E܋@;E�u�   ��    ����t�E��U܉P�E܋U��P�   �oM  �E���E؋E؋ �E܃}� u�E���E؋E؋ �E܃}� t�   ��    ��tg��EԉE؋E؋ �E܋E܃��EԋEԋ ��u�E܃��EԋEԋ ��t�   ��    ��u��E�@;E�������t�E��     ���L  �}� �E  �E�@��L��    �EЉE��E�� ;E�u9�E��U܉�E�� ������t\�E�P�E�@�   �������!E�P�9�E�@;E�������t!�E��@;E�u�E��U܉P��E��U܉P��,L  �}� ��   �E�@;E���������   �E܋U��P�E�@�E��}� ����t,�E�@;E�������t�E܋U��P�E��U܉P���K  �E�@�E��}� ����t,�E�@;E�������t�E܋U��P�E��U܉P��K  ��{K  �   ���P��   ��!�;E�v;�U��EЃ��E�P�U��EE�ЋM��UыU�ʋR���P�  �E���E�P�E����E��P�U��E�E���E�������   �E����E��E������    �EЃ��E��E��EЋE��E�����Ѓ���u�E��E��   �����	E��(�E��P�E�@9�������t�E��@�E���mJ  �E��U��P�EЋU��P�E��UЉP�E��U��P�  �E���|����E�����x�����x��� u	�E�    �R��x�����  v	�E�   �=�    ��x�����)Ѓ���t�����t���� ��t��������E����ЉE̋Ẽ�L��    �EЉ�p�����|����ỦP��|����@    ��|����P��|����P�E�P�Ẻ���Ѓ���u_�E�P�E̻   �����	E�P��p�����|������|�����p����P��|�����|����P��|����P��|����P�t  ��p���� �Eȃ}�t�    �E���)Ѓ�����    �E������EċEȋ@���;E���   �    ���Eĉ��������    �E�Љ�l����eċ�l���� ��t��l���� �E���   �E�@;�l���������t@��l�����|������|����UȉP��|�����|����P��|����P��|����P�   �)H  �Eȋ@��h����E�@;E�w�E�@;�h���w�   ��    ����tH��h�����|����P��h����P�EȉP��|�����h����P��|����UȉP��|����@    �
�G  ������   �E���
�G  �    �Ĕ   []�U��S��d�E�P�E�@��!ЉE���E؉EԋEԉEЋE�UЃ�L���E�E�E��E�@���+E�E��#�E�@���+E�E̋E�;E�s�ẺE�E�E��E�@��t�E�@��E�@�E�}� ����u��E�@;E���������  �U��EЉEȋE�;E���������  �E��@�EċE��@;E�tb�E��@�E��E��@�E�E�@;E�w�E��@;E�u�E�@;E�u�   ��    ����t�E��U�P�E�U��P�   �=F  �E����E�E� �E�}� u�E����E�E� �E�}� t�   ��    ��tg��E��E�E� �E�E���E��E�� ��u�E���E��E�� ��t�   ��    ��u��E�@;E�������t�E��     ��E  �}� �E  �E��@��L��    �EЉE��E�� ;E�u9�E��U��E�� ������t\�E�P�E��@�   �������!E�P�9�E�@;E�������t!�Eċ@;E�u�EċU�P��EċU�P���D  �}� ��   �E�@;E���������   �E�UĉP�E��@�E��}� ����t,�E�@;E�������t�E�U��P�E��U�P��D  �E��@�E��}� ����t,�E�@;E�������t�E�U��P�E��U�P��PD  ��ID  �   ���P��   ��!�;E�v;�U�EЃ��E��P�U�EE�ЋM�UыU�ʋR���P��   �E���E��P�E���EȉP�UȋE�E��E�@�E��}� ��   �E�@�E��E����E��E������    �EЃ��E��E��E܋E��E�����Ѓ���u�E��E��   �����	E��(�E��P�E�@9�������t�E��@�E���.C  �E��U��P�E܋U��P�E��U܉P�E��U��P�E�U�P�E�UȉP�   �E�����B  ��d[]�U��VS��p��[��u	�������t��|]����t#�   ��]��t��h�]蹿������u�   ��    ����  �������   ;E��  �   ���P��   ��!Ѓ���;Ev�   ���P��   ��!���E���   ЍP��   ��!ЉE��E����E��[�E����ЉE�E������   �E��������E�E�������[���E��E��@�E܋E܋@�E؋E�;E�u��[�E�   �������!У�[�A��[;E�w�E؋@;E�u�   ��    ����t�E؋U��P�E��U؉P��RA  �E������E܉P�E��    �E�ЋU��    �U�ʋR���P�   �E�ЉE��  ��[;E��@  �}� ��  �E�U����E�   ����؍ �E�   ��������	�!ЉEԋE���#EԉE���EЉE̋ẺEȋE�������[���EċEċ@�E��E��@�E��E�;E�u��[�EȻ   �������!У�[�A��[;E�w�E��@;E�u�   ��    ����t�E��UĉP�EċU��P��@  �E���+E��E��E����E��P�U��E�ЉE��E����E��P�U��E�E����[�E��}� ��   ��[�E��E����E��E�������[���E��E��E��[�E�����Ѓ���u��[�E��   �����	У�[�'�E��P��[9�������t�E��@�E���:?  �E��U��P�E�U��P�E��U�P�E��U��P�E���[�E���[�   �E�ЉE��
  ��[��t#���u�h�[�[������E�}� t�   ��    ��t��  �}�   ���P��   ��!�����;Ew	�E������V�E���   ЍP��   ��!ЉE��[��t#���u�h�[�-������E�}� t�   ��    ��t�Q  ��[;E���   ��[+E��E���[�E��   ���P��   ��!�;E�wH�U��E�У�[��[�E��E���[�E����E��P�U��E�E���E����E��P�C��[�E���[    ��[    �E����E��P�U��E�ЋM��U�ʋR���P�   �E�ЉE��}��[;E�v]��[+E��[��[�E���[�E��U��E�У�[��[�E��E����E��P�E����E��P�   �E�ЉE�����u�h�[�d������E��|]����t
�    ��]�E���    �e�[^]�U��S��   �} ��  �   �؉EЉE��|]����t#�   ��]��t��h�]葹������u�   ��    ���o  ��[;E�w�E�@����t�   ��    �����%  �E�@����E��U�E�ЉEċE�@�����  �E� �E��E�@����u�   �E��E���  �E��؉E�ЉE��E�E��E��E���[;E���������  ��[;E��_  �E�������   �E�@�E��E�@�E��E����E��E�������[��;E�t��[;E�w�E��@;E�u�   ��    ������   �E�;E�u��[�E��   �������!У�[�^�E�������[��;E�t��[;E�w�E��@;E�u�   ��    ����t�E��U��P�E��U��P�
�:  �:  �e  �E�E��E��@�E��E��@;E�ta�E��@�E��E��@�E��[;E�w�E��@;E�u�E�@;E�u�   ��    ����t�E��U�P�E�U��P�   �+:  �E����E�E� �E�}� u�E����E�E� �E�}� t�   ��    ��tf��E�E�E� �E�E���E�E� ��u�E���E�E� ��t�   ��    ��u���[;E�������t�E��     ��9  �}� �<  �E��@��L���[�E��E�� ;E�u8�E��U��E�� ������tZ��[�E��@�   �������!У�[�8��[;E�������t!�E��@;E�u�E��U�P��E��U�P���8  �}� ��   ��[;E���������   �E�U��P�E��@�E��}� ����t+��[;E�������t�E�U��P�E��U�P��8  �E��@�E��}� ����t+��[;E�������t�E�U��P�E��U�P��H8  ��A8  �G�Eċ@����u9�E��[�Eċ@����EĉP�E����E�P�U�E�E����  ���  �E�;E�s�Eċ@����t�   ��    ������  �Eċ@������  ��[;E�um��[�E�У�[��[�E��E���[�E����E�P��[;E�u��[    ��[    ��[;E�s��j h�[�������;  ��[;E�u@��[�E�У�[��[�E��E���[�E����E�P�U�E�E����  �Eċ@����E��E�E��E�������   �Eċ@�E��Eċ@�E��E����E��E�������[��;E�t��[;E�w�E��@;E�u�   ��    ������   �E�;E�u��[�E��   �������!У�[�^�E�������[��;E�t��[;E�w�E��@;E�u�   ��    ����t�E��U��P�E��U��P�
��5  ��5  ��  �Eĉ�|�����|����@��x�����|����@;�|���t|��|����@��t�����|����@�E��[;�t���w&��t����@;�|���u�E��@;�|���u�   ��    ����t��t����U��P�E���t����P�   �D5  ��|������E܋E܋ �E��}� u��|������E܋E܋ �E��}� t�   ��    ��tf��E؉E܋E܋ �E��E����E؋E؋ ��u�E����E؋E؋ ��t�   ��    ��u���[;E�������t�E��     ��4  ��x��� ��  ��|����@��L���[��p�����p���� ;�|���uA��p����U����p���� ������tl��[��|����@�   �������!У�[�G��[;�x���������t-��x����@;�|���u��x����U��P���x����U��P���3  �}� ��   ��[;E���������   �E���x����P��|����@��l�����l��� ����t4��[;�l���������t�E���l����P��l����U��P��^3  ��|����@��h�����h��� ����t4��[;�h���������t�E���h����P��h����U��P��3  ��3  �E����E�P�U�E�E����[;E�u�E��[��  �,�Eċ@����EĉP�E����E�P�U�E�E���E�������   �E�����d�����d���������[����`�����`����Eԋ�[��d�������Ѓ���u ��[��d����   �����	У�[�-��`����P��[9�������t��`����@�E��� 2  ��`����U�P�EԋU�P�E�UԉP�E�`����P��  �E�\����E�����X�����X��� u	�E�    �R��X�����  v	�E�   �=�    ��X�����)Ѓ���T�����T���� ��T��������E����ЉEЋEЃ�L���[��P�����\����UЉP��\����@    ��\����P��\����P��[�EЉ���Ѓ���u^��[�Eл   �����	У�[��P�����\������\�����P����P��\�����\����P��\����P��\����P�q  ��P���� �Ẽ}�t�    �E���)Ѓ�����    �E������EȋE̋@���;E���   �    ���Eȉ��������    �E�Љ�L����eȋ�L���� ��t��L���� �E���   ��[;�L���������t@��L�����\������\����ỦP��\�����\����P��\����P��\����P�   �/  �E̋@��H�����[;E�w��[;�H���w�   ��    ����tH��H�����\����P��H����P�ẺP��\�����H����P��\����ỦP��\����@    �
�9/  �������[����[��[������t��h�[�`�������/  �|]����t
�    ��]�]���U����E�    �} t/�E�E�E�EEf�  ��t�E��    �u;Et�E��������u��������E��}� t+�   �؉E�Ћ@����t���u�j �u��4  ���E���U��S��   �E�    �E�@����E�U�E�ЉE��E�@;Ew*�E�@����t�E;E�s�E��@����t�   ��    �����;  �E�@����u�u�u�u�u�������E��  �E�;E��   �E�+E�Eܸ   ���P��   ��!�;E�w�U�EЉE؋E�@��E���E�P�U�EЋM�UʋR���P�E؋@��E܃��E؉P�U؋E�ЋM؋U�ʋR���P���u��u��u�������E�E��X  �E�@;E���   �E�P�E��;Evx�E�P�E�ЉEԋE�+E�EЋU�EЉE̋E�@��E���E�P�U�EЋM�UʋR���P�EЃ��ẺP�E�ỦP�E�UЉP�E�E��  �E�@;E��%  �E�@�EȋU�E��;E�  �U�E��+E�Eĸ   ���P��   ��!�;E���   �U�EЉE��U��E�ЉE��E�@��E���E�P�U�EЋM�UʋR���P�Eă��E��P�U��E�Eĉ�E��@����E��P�E�UĉP�E�U��P�O�U�E�ЉE��E�@��E����E�P�U�E�ЋM�U�ʋR���P�E�@    �E�@    �E�E��  �E��@�����w  �E��@����E��U�E��;E�Z  �U�E��+E�E��E�������   �E��@�E��E��@�E��E����E��E������    �EЃ�;E�t�E�@;E�w�E��@;E�u�   ��    ������   �E�;E�u�E��E��   �������!E��c�E������    �EЃ�;E�t�E�@;E�w�E��@;E�u�   ��    ����t�E��U��P�E��U��P�
�*  �*  �p  �E��E��E��@�E��E��@;E�tb�E��@�E��E��@�E��E�@;E�w�E��@;E�u�E��@;E�u�   ��    ����t�E��U��P�E��U��P�   �)  �E����E�E� �E��}� u�E����E�E� �E��}� t�   ��    ��tg��E�E�E� �E��E����E�E� ��u�E����E�E� ��t�   ��    ��u��E�@;E�������t�E��     ���(  �}� �E  �E��@��L��    �EЉE��E�� ;E�u9�E��U���E�� ������t\�E�P�E��@�   �������!E�P�9�E�@;E�������t!�E��@;E�u�E��U��P��E��U��P��D(  �}� ��   �E�@;E���������   �E��U��P�E��@�E��}� ����t,�E�@;E�������t�E��U��P�E��U��P���'  �E��@�E��}� ����t,�E�@;E�������t�E��U��P�E��U��P��'  ��'  �   ���P��   ��!�;E�v=�U�E�ЉE��E�@��E����E�P�U�E�ЋM�U�ʋR���P��U�EЉE��E�@��E���E�P�U�EЋM�UʋR���P�E��@��E����E��P�U��E�ЋM��U�ʋR���P���u��u��u��������E�E���&  �E�]���U���H�E�    �   ���P��   ��!�;Ev�   ���P��   ��!ЉE�E��#E��t�   ��E���e��E�;Er��E��E�   ���P��   ��!�����+E;Ew"�} �*  e�    ������2   �  �   ���P��   ��!Ѓ���;Ev�   ���P��   ��!���E���   ЍP��   ��!ЉE�U�E¸   ���H��   ��!�Ѓ��E���u��������E�}� ��  �   �؉E�ЉE�E���  ����t3�E���  �   ���t�E�  ��P�D�������t�   ��    ��t
�    �  �E�P��E�!Ѕ��  �E�P��E�ЉE��!к   )ЉE��U��E�)Љ��   ���P��   ��!�9�s
�U��E���E��E܋E܉E؋U܋E�)ЉEԋE�@���+EԉEЋE�@����u�E��E�E؉�E؋UЉP�t�E؋@��EЃ��E؉P�U؋E�ЋM؋U�ʋR���P�E�@��Eԃ��E�P�U�E�ЋM�U�ʋR���P���u��u��u��������E؉E�E�@������   �E�@����E̸   ���P��   ��!E��;E���   �E�+E�EȋU�E�ЉEċE�@��E���E�P�U�E�ЋM�U�ʋR���P�Eċ@��Eȃ��EĉP�UċE�ЋMċU�ʋR���P���u��u��u�������   �E�ЉE�E���  ����t�E�  �    ��E���U���8��[��u	������t��} t�} u�E�  �E�E��E�    �|�} u��j �������  �E�    �E��    �   ���H��   ��!ȃ���9�s�   ���P��   ��!���E�����   ЍP��   ��!ЉE�E����tf�E� �   ���J��   ��!ʃ���9�s�   ���P��   ��!���E� ���   ЍP��   ��!ЉE�E�E�E��   �E�    �E�    �E�    �s�E؍�    �EЋ �   ���J��   ��!ʃ���9�s�   ���P��   ��!��'�E؍�    �EЋ ���   ЍP��   ��!�E��E��E�;Eu��U��E�ЉE��E�    �E܃���P�,������EЃ}� t�E���  �E���  �}� u
�    ��  �E���  ����t3�E���  �   ���t�E�  ��P�ŝ������t�   ��    ��t
�    �  �   �؉E�ЉE�E�@����E�E����t�E��+E��Pj �u��n&  ���}� u5�U�E�ЉE̋E�+E��EȺ   �E�ЉE��Eȃ��ẺP�E��E��E�    �E؍�    �E�й   �U�ʉ�E��;E���   �}� t�E�E��o�E؍�    �EЋ �   ���J��   ��!ʃ���9�s�   ���P��   ��!��'�E؍�    �EЋ ���   ЍP��   ��!ЉE܋E�)E�E܃��E�P�E�E��!�E���E�P��E���  ����t�	�E������E�  �    ��E���U���8�E�    �E���  ����t,�E���  �   ���t�E�  ��P�ޛ������u�   ��    ���{  �E��    �EЉE�E�E��  �E� �E�}� ��   �   �؉E�ЉE�E�@����E��E��     �E�@;E�w�E�@����t�   ��    ������   �E���E܋E�@����E�ЉE؋E�;E�th�E܋ �   �U��9�uU�E؋@����E�ЉEԋE�@��Eԃ��E�P�U�E�ЋM�U�ʋR���P�   �E�E܉�����u��u��u��������|  �E��E�;E�������E�P�E�@9�v��j �u�������E���  ����t�E�  �    ��E���U���(�E�    �} u���u�)������E��  �   ���P��   ��!�����;Ewe�    ������2   �u  �   ���P��   ��!Ѓ���;Ev�   ���P��   ��!���E���   ЍP��   ��!ЉE�   �؉EЉE��E��[�E苀�  ����t,�E荐�  �   ���t�E��  ��P�F�������u�   ��    ����   j�u��u��u��������E�E苀�  ����t�E��  �    ��}� t�   �E�ЉE��r���u��������E�}� t[�E�@����E�@����u�   ��   )ЉE��E�;Es�E���E��P�u�u��   �����u�������E���U���(�E�    �} �.  �   ���P��   ��!�����;Ewe�    ������2   ��   �   ���P��   ��!Ѓ���;Ev�   ���P��   ��!���E���   ЍP��   ��!ЉE�   �؉EЉE��E��[�E苀�  ����t,�E荐�  �   ���t�E��  ��P��������u�   ��    ��tCj �u��u��u���������E�E苀�  ����t�E��  �    ��E�;E�u�E�E�E���U����   ;Er���u�	���������u�uh�[�)�������U����E�    �   ;Eu���u��������E��   �E���E��E���E�}� u�}� t�E���#E���t
�   �   �   ���P��   ��!�����+E;ErI�   ���P��   ��!�;Ev�   ���P��   ��!ЉE���u�uh�[�^������E�}� u�2   ��E�U��    ��U�����[��u	������t���[�E���u�u���������U�����[��u	豖����t���[�E�U�E�ЍP��E���!Ѓ�P�u��m�������U����E�E���uj�E�P�uh�[�`����� ��U������uj �u�uh�[�=����� ��U������u�uh�[��������U����E�    ��[��u	�������t��|]����t#�   ��]��t��h�]�Ք������u�   ��    ��t,���uh�[�P������E��|]����t
�    ��]�E���U��p]]�U��t]]�U����x]�E��}� t�E���������U����} u��[��[��!ЉE��}�u	�E�    ���[�EЍP���[��!ЉE��E��x]�x]��U����E��h�[P�x������E�� U�����h�[�ۘ������U������u�u谕������U����} tI�   �؉EЉE��E��@����t*�E��@����E��@����u�   ��   )���    ��U�����F  �    ��U����} u�}u�E�����u�u��D  ����U������u�(   ���E�}� t���������u�
������    ��U����E����P�cB  �����u�   ���E�E�@ �E���U������u�  ���E�@0���u�Ѓ�������t������Z�E�@L%   ��t&�E�@��t�E�@L��y�E�@��P�d�������jXj �u�8  �����u�  ���    ��U�����jjX�������E�}� ue�    ������2   �    �(���u��u�u�   ���������t�    ��E���U������u�  ���E�}��u
������   �E�U��U�E�PL�E�@�E�@0���E�@  ��E�@$
��E�@(ŵ�E�@,��E�@8
��E�@4?��E�@@��E�@<ʴ���u��  ���    ��U����} u6�E�    ��]�E�����u��������	E�E��@T�E��}� u��E��-�E����P�Q@  �����u�   ���E�E�@ �E���U����E�@L%    ��t���u�  �����u�   ��    ��t������>�E�@L%   @��t���u�&   �����u�   ��    ��t�������    ��U��S��$�E�@L%   @��u
�    �E  �E�@L����u0e�    ������   �E�@L   �E�PL������  �E�@$��u0e�    ������   �E�@L   �E�PL�������   �E�    �E�@�E��E�    �   �E�@$�U�+U��M�Y�M�ك��uRQ�Ѓ��E��U�E�E���u�E�@L   �E�PL�E������B�E����E����	Ѕ�u�E�@L   �E�PL�E�������E�E��E�;E��n����E�@L%�����E�PL�E�@    �E�]���U��E� ]�U�����jjX�������E�}� ue�    ������2   �    �5���u��u�u�&   ���E��}� u���u��f������    ��E���U������u�	  ���E�}��u�    �V���u��u�@  ���E��}��u�    �5���u�u�u��)�����������t�E����u��  ���    ��U����E�E��E���P�u�u��  ���E�E���U����E����P�=  �����u�u�   ���E�E�@ �E���U��S���E�E��E�@L%   ��u"���u�	  ���������t
������  �E�@<u3�ujj�E�P�>  ��������t
�������   �E�����   �E�@L%    ��t"���u�[  ���������t
������   �E�P�E�@9�u���u�x������������t������j�E�@L   @�E�PL�E�X�E�@�H�U�J��E���E�@<u'�E�<
u���u�������������t�������E����]���U������u��  ���E��uj�u��u��  ���E��E�;E�u�E���������U����E����P�Q;  ���u�u�u�u�   ���E�E�@ �E���U���8�} t�} u
�    �+  �E�@L����u0e�    ������   �E�@L   �E�PL�������  �E�@L%   ��u"���u�  ���������t
������  �E�@<�C  �E�@L%   @��t"���u��������������t
������}  �E�@ ��u0e�    ������   �E�@L   �E�PL������C  �E�@L    �E�PL�E�@L%�����E�PL�E�    �E�E�E��E�    ��E�@ �M�U�ʃ��u�u�R�Ѓ��E؉U܋E�E؅�u�E�@L   �E�PL�E������B�E܃���E؃��	Ѕ�u�E�@L   �E�PL�E�������E�E�E�;E��u����E��    �u�k�E�E��E�    �Q�E��E�E��E�    �2���u�  ���Ẽ}��u�E��-�UЋE�E�ЋÜ�E��E�;ErƃE��E�;Er��E��U����E��uRP�u�   ����U���(�E�E��E�E�E����P�8  ���u�u��u��u�   ���E�E�@ �E���U���(�E�E��E�E�E�@(��t�E�@(�u�u��u��u�Ѓ��E��e�    ������>   �E������E���U������u�   ����U����E����P��7  �����u�   ���E�E�@ �E����U����E�@,��t�E�@,���u�Ѓ��E��e�    ������>   �E������E����U����E����P�7  ���u�u�u�u�   ���E�E�@ �E���U���(�} t�} u
�    �,  �E�@L����u0e�    ������   �E�@L   �E�PL�������  �E�@L%   ��u"���u�  ���������t
������  �E�@<�A  �E�@L%    ��t"���u�  ���������t
������~  �E�@$��u0e�    ������   �E�@L   �E�PL������D  �E�@L   @�E�PL�E�@L%�����E�PL�E�E�E��E�    �   �E�@$�M�U�ʃ��u�u�R�Ѓ��E��U�E�E���u�E�@L   �E�PL������   �E����E����	Ѕ�u�E�@L   �E�PL������   �E�E�E�;E��s����E��    �u�n�E�E��E�    �T�E��E�E��E�    �5�U؋E�E��� �����uP�N������������t�E���E��E�;ErÃE��E�;Er��E��U����E����P��4  �����u�b  ���E�E�@ �E���U����   ��]�U�PP��]�E�PT�E��]�s   ��U����N   ��]9Eu�E�@T��]�E�@P��t�E�@P�U�RT�PT�E�@T��t�E�@T�U�RP�PP�   ��U�����h�]�?4  ����U����] ]�U����E�    �E� ����rt��wt��at��E�   �,�E�R   �#�E�b   �e�    ������   ������d�L�E� ����bt��tt��+u�M��.�e���M��$�e���M��e�    ������   �������E�E� ������u��E���U����E����P�W3  �����u�u�T������E�E�@ �E���U���h    jj �u�y   ��������t�    �)h    jj �u�U   ��������t�    ��������U����E����P��2  ���u�u�u�u�   ���E�E�@ �E���U����E�@<t&�E�@��t�E�@L��y�E�@��P��������} uO�} u	�E    ��}w�E�   ���u�������E�} u������{�E�@L   ��E�PL��E�@L%����E�PL�E�U�P�E�E�P�E�U�P�E�@    �E�@    �E�@    �E�@L   �E�PL�    ��U����E�E��E���P�u�u��  ���E�E���U�����h��	�|������j �2  ����U�����D��jXj P�
  ����D��Phh�	j ���������Dh   jh@^P�9�������D��jXj P�q
  ����D��Phj�	j��������Dh   jh�bP���������D��jXj P�*
  ����D��Phj�	j�T�������Dh   jh@gP��������U�����]�E��M�E�@T�E��E�����P�0  ��������t#���u����������u���������E��@ �E��E�}� u���U����E� ��P�;  ����U��E�@L%   ��t�   ��    ]�U��E�@L%   ��t�   ��    ]�U������u�n�������U����E� ���u�uP��  ����U����} uF���u�M������E�}��u�    �Z�E�@Lf�  �E�PL�E�PL�E�	E�PL�E�2���u��������E��}� t�    ����u�u�u�B�������U����E�E��E�E�E� �u�u��u�P�n
  ����U����E� ��P��  �����U����E� ���u�uP��  ����U����E����P�.  �����u�u�  ���E�E�@ �E���U����E����P�[.  �����u�u�u�2   ���E�E�@ �E���U����u�uj�u��������    ��U����E�@L����u-e�    ������   �E�@L   �E�PL�������u�uh���u��  ����U����E�E�E�P�E�@9�sV�E�P�E�@)ЉE��E;E�s�E��E��E�E��E�@Ѓ��u��uP��  ���E�P�E�E�P�E�P�EE�P�E�    ��U���(�E�E�} t�E����    �E��E�    �E�    �u�uh��E�P�!  ���E�} t�U�E���  �E���U����u�uj��u��������U�����j��R-  ����U�����|����0  ���u�2-  ��U�����h   �ټ�����E����u��C-  �����u��y
  ���E��E�    ���u��  ���E�}��  w&�E����P脼�����E���u��u��.  �����u��������E���U���H��h   �G������Eȃ}� u
������K  ���u��",  ���EȉE��E�   �   ��E��E�� ��t�E�� ����P�Vz������u��E� �E� �q�E�� <"u�E����t
�u��E� �N�E�� <\u�E����t�E��3�E�� ����P��y������t�E����t�E����u�E� �E��E�� ��u��E��E�� ���@����E�������P�?������Eă}� u
������C  �8����Eĉ�EȉE��E�   ��   ��E��E�� ��t�E�� ����P�Py������uًE�P�U��    �E�E��E� �E� �q�E�� <"u�E����t
�u��E� �N�E�� <\u�E����t�E��3�E�� ����P��x������t�E����t�E����u�E� �E��E�� ��u��E�� ��u��E�P�U��  �E�� �������E��    �E���     �E�   ��   �E���    �E�Ћ �E����u���  ���E��E� �E�    �   �Eۃ���tI�UԋE��� <\u:�EԉE���UЋE�EЍH�E��� ��E��E�;E�r܃m��m��E��X�Eۃ���tI�UԋE��� <"u:�EԉE���ŰE�E̍H�E��� ��E��E�;E�r܃m��m��E� ��E� �E��E�;E��D����E��E�;E�������E�U���E�Uĉ�    ��U�����h �	�s������j �)  �����	�����	��U�����h��	��r������j ��(  ���L�	���L�	��U����E�E���E�� �U8�u�E���E��E�P��U������uظ    ��U����E�E��E�E��E�    �F�U��E����M�E��� 8�v�   �2�U��E����M�E��� 8�s�������E��E�;Er��    ��U����E�E��E�E���E��P�U��U��J�M����E�P��U������u׋E��U����E;EvI�E�P��EЉE��E�P��EЉE���E��P��U��U��J��M����E�P��U������u��7�E�E�E�E���E��P�U��U�J�M����E�P��U������u׋E��U����E�E���U��EЋU��E�P��U������u�E��U����E�E��E�E��E�� �E��E�� �E��}� u�}� u�    �*�E�:E�s�������E�:E�v�   �
�E��E����U�����h��	�p������j �&  ����U����E�P�U�U�J�M���E� ��uߋE�  �E]�U��(�	]�U����E�    ��E��U�E��� ��u�E���U������u�u�u�$  �����u��������U������u�uhн	��  ���    ��U������uh��	�  �����u�u�*��������u�W�������U�����%  �E��U�U��E��E���U������u�H%  ���E�}� u�    �3�}�ue�    ������   �e�    ������   �������U���8�E�EЋE�Eԃ}u	�E�    ��}u	�E�   ��}u�E�   ���E�P�u��u��u��u��&  �� �E�U�E��u�E�U��:�E��ue�    ������   �e�    ������   ������������U����E�    ���M�QRP�u�u�%  �� �E�E���u�E���W�E���ue�    ������   �0�E���ue�    ������   �e�    ������   ������������U������E�P�u�%  ��������t�E��e�    ������2   �������U������u�&  ����U����E�    ���M�QRP�u�u�_&  �� �E�E���u�E���W�E���ue�    ������   �0�E���ue�    ������   �e�    ������   ������������U����E�    �E��@��t�E�E�E�P�U� �E���E�P�u�u�|#  ���E��E��u�E��5�E��ue�    ������.   �e�    ������   �������U����} u�@k.�Ak �@k�   ���u�������E��}� u�@k.�Ak �@k�o�E��P��EЉE��
�E��  �m��E�;Er
�E�� </t�E� ��u�@k/�Ak �@k�$��j/�u��   ���E�}� u�E��E����U��]�U�����j �a���U��S��$�E�@L%    ��u
�    �P  �E�@L����u0e�    ������   �E�@L   �E�PL������  e�    �������E��E������E������E�@(��t�E�@(jj j �u�Ѓ���E��U�e�    ������M��E�    �}� ��   �E�P�E�@)ЉE�E��U�M�    9�r9�w9�r�M�    �E��U�)���
�    �    �E؉U܋E�@(j�u��u��u�Ѓ�����t�E�@L   �E�PL�E�@    �E�@    �E�@L%���߉E�PL�E�]���U��S��$�E�@L%   ��u"���u�7������������t
������b  �E�@<u3�ujj�E�P������������t
������0  �E����$  �E�@L%   @��t"���u�J������������t
�������   �E�@L    �E�PL�E�P�E�@9���   �E�   �E�@;E�w�E�    �E�@ �U�R+U�M�Y�M�ك��uRQ�Ѓ��E�U�E�E��u�E�@L   �E�PL������b�E����E���	Ѕ�u�E�@L   �E�PL������4�U�E�E�P�E�U�P�E�X�E�@�H�U�J�� ���]���U��S���E�@L%   ��u"���u�������������t
������>  �E�@<u0e�    ������   �E�@L   �E�PL������  �E�@L%   @��t"���u�������������t
�������   �E�@L    �E�PL�E�@L%�����E�PL�}�u
������   �E�E��E�@��ue�E�P�E�@)ЉE��E�@+E��E�}� u������`�U��E�@�M�Y�M�ك�RPQ�������E�U�P�U�E�E�P�E�P�E�@�H��E�H�E�@��E���E��]���U����E�E�E��P�u�   ����U������u�������E�E����E����u�葬�����E��u�u�u��u�����������u��f�������u��|�������U����E�    �E� �E��#�U��������E�� ����0ЉE��E��E�� </~
�E�� <9~ɋE�U���E���U��S��4�E�EЋE�EԋE�EȋE�E��E�   �EЋUԉE�U���u��u��u��u��#�����E�U�E��E�U�;U�w�;U�r;E�s͋E�E��L�E�P��E��EЋU��u��u�RP�$�����E�� ��u��u��u��u��%#�����EЉUԃm��}� u��E�]���U��WVS��,  �E��$����E�    ��  ��$���� <%�`  ��$�������$�����$���� ������t�E���  ��$���� <%��   ��$�����jP�u�E�Ѓ��ǃ��������Ѐ� ��������������������	�������t
������a  �E���$�������$�����$���� ������t�E��4  �  �E� �E� �E� �E� �E� �E� ��$���� ���� ��w:��x�	���E��E��'�E��E���E��E���E��E��	�E��E���}� t)��$�������$�����$���� ������t�E��  �}� �u����E�    ��$���� <*u7�U�B�E��E؋�$�������$�����$���� ������t7�E��E  ��$���� </~"��$���� <9����$���P��������E��E�   �E� ��$���� <.��   ��$�������$�����$���� ������t�E���  �E���$���� <*u7�U�B�E��Eԋ�$�������$�����$���� ������t7�E��  ��$���� </~"��$���� <9����$���P�������E��E�    ��$���� <huv��$�������$�����$���� ������t�E��  ��$���� <hu4�E�   ��$�������$�����$���� ��������  �E���  �E�   �  ��$���� <luv��$�������$�����$���� ������t�E��  ��$���� <lu4�E�   ��$�������$�����$���� �������  �E��Y  �E�   ��   ��$���� <ju5��$�������$�����$���� ������t�E��  �E�   �   ��$���� <zu2��$�������$�����$���� ������t�E���  �E�   �|��$���� <tu2��$�������$�����$���� ������t�E��  �E�   �=��$���� <Lu0��$�������$�����$���� ������t�E��W  �E�   ��$���� �Eˋ�$���� ����A��7��  ����	���}�dt
�}�i��   �E��}���   �E�����	� ���U�B�E���E��U��   �U�B�E�����E��U��   �U�B�E����E��U��   �U�B�E���E��U��t�U�B�E��R�E��U��^�U�B�E��R�E��U��H�U�B�E��E��E�    �1�U�B�E���E��U��e�    ������   ������%  ��   �E� �}���   �E�����	� ���U�B�E��E��E�    ��   �U�B�E����E��E�    �   �U�B�E����E��E�    �   �U�B�E��E��E�    �t�U�B�E��R�E��U��^�U�B�E��R�E��U��H�U�B�E��E��E�    �1�U�B�E���E��U��e�    ������   ������$  �}� t�E��Uą�y�   ��    ��W����}�pu�E�x�E��}�xu�E�   �E�0�	�:�}�Xu�E�   �E�A�	�$�}�ou�E�   �E�R�	��E�
   �E�\�	�E���������W��� t�E��U��؃� ����E��Uă��u�SQRP�����P������ ��H���ǅL���    �E�    �}� u�}� u	��W��� t�E��}� t�}�xt�}�Xu�E��}� t
�}�ou�E��E؉Ɖ����E���������H�����L�����9�9�|9�s��H����E�ЉE��E������   �E߃�����   �E�    �V��jhg�	�u�E�Ѓ��ǃ��������Ѐ� ��������������������	�������t
������Z  �E��E��E��Ɖ����Eؙ+�H����L������ӋE��)�Ӊȉ�9��x���9�9��l�����W��� tW��jhi�	�u�E�Ѓ��ǃ��������Ѐ� ��������������������	�������t
������  �E��   �}� tT��jhk�	�u�E�Ѓ��ǃ��������Ѐ� ��������������������	�������t
������`  �E��X�}� tR��jhg�	�u�E�Ѓ��ǃ��������Ѐ� ��������������������	�������t
������  �E��E������   �}� ��   �E�    �V��jhm�	�u�E�Ѓ��ǃ��������Ѐ� ��������������������	�������t
������  �E��E��E��Ɖ����Eؙ+�H����L������ӋE��)�Ӊȉ�9��x���9�9��l����}� �
  �}�xt
�}�X��   ��jhm�	�u�E�Ѓ��ǃ��������Ѐ� ��������������������	�������t
�������  �E��}�xuN��jho�	�u�E�Ѓ��ǃ��������Ѐ� ��������������������	�������tX������  ��jhq�	�u�E�Ѓ��ǃ��������Ѐ� ��������������������	�������t
������>  �E��^�}� tX�}�ouR��jhm�	�u�E�Ѓ��ǃ��������Ѐ� ��������������������	؅�����t
�������  �E���H�����P�����P�u�E�Ѓ���3�H�����x�����3�L�����|�����x�����|�����	؅�����t
������  ��H����E�ЉE�}� ��   �E�    �V��jhg�	�u�E�Ѓ��ǃ���p����Ѐ� ��t�����p�����t�����	؅�����t
������  �E��E��E��Ɖ����Eؙ+�H����L������ӋE��)�Ӊȉ�9��x���9�9��l����8  �E̅�t��t�,�U�B�E��}��9�U�B�E��J�R�E��U��M��e�    ������   ������n  �m�����������G�����G��� t�m����}��m��-p�	������s-�m�ٽ�����������f������٭����߽8���٭�����k�m��-p�	��ٽ�����������f������٭����߽8���٭������8����� ��h�����<���5   ���l�����h�����l�����8�����<�����8�����<�����8�����<����m�٭����߽����٭����߭�����m����]�����E����	���]��E�٭����߽����٭����߭����ݝ����݅�����E�������z�������u��E����	������s�E�٭����߽0���٭�����U�E����	��٭����߽0���٭������0����� ��`�����4���5   ���d�����`�����d�����0�����4�����0�����4�����0�����4�����h\�	j j
��<�����8��������P�|����� ��,�����h\�	j j
��4�����0���������P�O����� �E��E�;E�s�EԉE��E�    �}� u�}� u	��G��� t�E��}� t�E��-�E�    ��������E��� <0t�E���E��E�;E�r܋M؋U���,���E��9�s�U���,���E�ЉE��E������   �E߃���t}�E�    �V��jhg�	�u�E�Ѓ��ǃ���X����Ѐ� ��\�����X�����\�����	�������t
������-	  �E��E��M��E�+�,����E�)E�)�9�r���G��� tW��jhi�	�u�E�Ѓ��ǃ���P����Ѐ� ��T�����P�����T�����	؅�����t
������  �E��   �}� tT��jhk�	�u�E�Ѓ��ǃ���H����Ѐ� ��L�����H�����L�����	�������t
������S  �E��X�}� tR��jhg�	�u�E�Ѓ��ƃ���@����Ѐ� ��D�����@�����D�����	؅�����t
�������  �E��E������   �E߃�����   ǅ|���    �Y��jhm�	�u�E�Ѓ�������8����Ѐ� ��<�����8�����<�����	�������t
������}  �E���|�����|����E�+�,����E�)E�)�9�r�����,��������P�u�E�Ѓ����Ӌ�,����    ��1ǉ�0���1Ӊ�4�����0�����4�����	؅�����t
�������  �U䋅,���ЉE�}� u��4����0������8  ��jhs�	�u�E�Ѓ��ƃ���(����Ѐ� ��,�����(�����,�����	�������t
������|  �E����u�������P�u�E�Ѓ����ӋE��    ��1ǉ� �����1щ�$����� �����$�����	؅�����t
������  �U�E�ЉE�ǅx���    �Y��jhm�	�u�E�Ѓ��Ã�������Ѐ� �����������������	�������t
������  �E���x����}� t�E�+E���   ;�x���w��}� ��   ǅt���    �Y��jhg�	�u�E�Ѓ��ƃ�������Ѐ� �����������������	؅�����t
������.  �E���t�����t����E�+�,����E�)E�)�9�r��p  �E̅�t��t�&�U�B�E��������0�U�B�E��������e�    ������   ������  �E����tsǅp���    �Y��jhg�	�u�E�Ѓ�����������Ѐ� �����������������	�������t
������G  �E���p����E؃�;�p������j������P�u�E�Ѓ��Ã��� ����Ѐ� ������� ����������	؅�����t
�������  �E��}� tsǅl���    �Y��jhg�	�u�E�Ѓ��ǃ��������Ѐ� ��������������������	�������t
������z  �E���l����E؃�;�l�����"  �E̅�t��t�&�U�B�E���h����0�U�B�E���h����e�    ������   ������  ����h�����������d����E�;�d���s	��d����E��E����txǅ`���    �Y��jhg�	�u�E�Ѓ��ƃ��������Ѐ� ��������������������	؅�����t
������{  �E���`�����`����E�+�d���9�r��}� t�E�;�d���s	�Eԉ�d�������d�����h����u�E�Ѓ����Ӌ�d����    ��1ǉ�������1щ�������������������	�������t
�������  �U䋅d���ЉE�}� ��   �E�;�d���vxǅ\���    �Y��jhg�	�u�E�Ѓ��Ã��������Ѐ� ��������������������	؅�����t
������f  �E���\�����\����E�+�d���9�r��}� txǅX���    �Y��jhg�	�u�E�Ѓ��ƃ��������Ѐ� ��������������������	�������t
�������   �E���X�����X����E�+�d���9�r��;�U�B�E���(�����(����E��e�    ������   ������   �Q��$�����jP�u�E�Ѓ������������Ѐ� ��������������������	؅�����t������>�E���$�������$�����$���� ������t�E����$���� �������E�e�[^_]�U����E�    ��U�E�M�E��� ��E��E�;Es�U�E��� ��u���U�E���  �E��E�;Er�E��U������u�������EЉE�E�� ��;Eu�E���E;E�u��    ��m�����U���j jj �u�M������U���j j�u�u� M������U���jjj �u��L������U���jj�u�u��L������U����E�E�E��Ph  �tL������U����E�E��E���Ph  �RL�����E���U����E�E�E��Ph  �-L����U�����j h  �L����U����E�E�E��Ph  ��K������U����E���Ph  ��K�����E��U���U���j j j �u�:   ����U���j j �u�u�    ����U����uj �u�u�   ����U���(�E�E�E�E�E�E�E��Ph  �WK�����} t�U��E��E���U����E�E��E�E��j �u��u��u�u�   �� ��U���8�E�EЋE�EԋE�E܋E�E��EЋUԉE�U�E܃�Ph  ��J�����} t�U�E��E��U���U���(�E�E�E�E븐0�E�E��Ph  �J�����E���U����E�E�E��Ph  �pJ�����E�E��E���U����E�E��E�E��j �u�u��u��u�   �� ��U���8�E�EЋE�EԋE�E܋EЋUԉE��U�E�E�E܃�Ph
  ��I�����} t�U�E��E��U���U�����j �u�   ����U����E�E�E��Ph  �I�����} t�U�E��E��U���U����E�E��E�E��j �u��u��u�u�   �� ��U���8�E�EЋE�EԋE�E܋E�E��EЋUԉE�U�E܃�Ph  �&I�����} t�U�E��E��U���U�����j h  ��H������f�f�f�f�f��U��S�(D���(D���t�v ��'    ���Ћ���u��[]�U���F���]�                                                                                ��������                                                                                                                                                                                                                                                                             ps2driver failed to register as    failed to allocate transfer memory area mouse did not ack set-default-settings command  mouse did not ack enable-mouse command                                          ��������                                                                                                                                                                                                                                                                             registering irq handlers                                           ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                             /var/log/ log.sys  [ ]                                             ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                           ��������                                                                                                                                                                                                                                                                             �� �P�����`�`�`�`� ������So  �	 �       �	���    L�`�                               ���М����������� �                        N9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE   	��,	                                                                ��`���`1p1@�p�0��1���������� �POSIX basic_string::erase %.*Lf %m/%d/%y %H:%M %H:%M:%S %s: __pos (which is %zu) > this->size() (which is %zu)   7 7�6�4@7@? ?�>�<`?�} }`|@|�u�u�u|�{�u�u�u�{�u�u�u�u�{p{P{�u�u�u@{`|py�u�u�u�u�u�u yx x�w0w�u�ux�u�u�u�u�v@v�u�u�u�u�u v�u�u�u�u`|P� ������� �Вp�@����	��St10ctype_base  �	�St9time_base    �	�St10money_base  �	4�St13messages_base   �	P�St12codecvt_base St7collateIcE  	a��
	St14collate_bynameIcE   	|�p�St8numpunctIcE  	���
	St15numpunct_bynameIcE  	����St7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE   	���
	                        St7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE   	@��
	St17__timepunct_cacheIcE    	���
	St11__timepunctIcE  	���
	St10moneypunctIcLb1EE                           �	��       �
	   �   St10moneypunctIcLb0EE           �	 �       �
	   �   St8messagesIcE                  �	`�       �
	   ,�   St23__codecvt_abstract_baseIcc9mbstate_tE                       �	��       �
	   H�   St14codecvt_bynameIcc9mbstate_tE    	 ��	St17moneypunct_bynameIcLb0EE    	0�@�St17moneypunct_bynameIcLb1EE    	\� �                        St9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE 	���
	                        St9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE 	 ��
	                        St8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE  	`��
	                        St15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE  	����                St8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE      �	 �       �
	   ��   St15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE  	��`�St15messages_bynameIcE  	����St18__moneypunct_cacheIcLb0EE   	���
	St18__moneypunct_cacheIcLb1EE   	 ��
	St16__numpunct_cacheIcE 	L��
	St21__ctype_abstract_baseIcE                    �	p�       �
	   ��       p�p�p���� �        ��0������ �        ��P�������@�p���                                ����0�����@�p���                                �P�`�`�����0�����P����`���        |�`���K N`Q�VPZ@a`d�Q    ��p���    ���� �                     �@G�G� ��������0�@�`�                @��G H�������� �P�������        �������`��                ��        ��������������                        $�@�P�@C`CpC�C�C�C�C                        P���P��������� �P�������                |������ ��������0�@�`�        ��0�����Н    <�@����B`D    ������)        ����)                `���@���@`�m0o                             ����p���@`�m0o     ��0�@���`��        ����    @�@�0�    d����                                            ��        ������������������������  St5ctypeIcE                 �	D	       �
	   ��       `	p��������0���������                             @       N9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEE    	�	�	                                    	����] H�Z�\ I�H P�K 30I�J�X                     "   7   Y   �   �   y  b  �  =  
  U  m  �*  /E  �o   �  % 1� B� s� �� (� ݊ =! ��5 �W �̌ ��� y�p)pT���~m��	8����ݥ�)�?�C_�sm�$�        St15basic_stringbufIcSt11char_traitsIcESaIcEE   	@	,	    St19basic_istringstreamIcSt11char_traitsIcESaIcEE   	�	�	St19basic_ostringstreamIcSt11char_traitsIcESaIcEE   	�	�St18basic_stringstreamIcSt11char_traitsIcESaIcEE    	 	�	    p	P���`1� p	�1`�@3�� 3��`200       �	        ���������	        �	�	�	�	        0       �	�������������	0�p�                        ,       �        ���������        L		 	`	        ,       �	�P����������	����                        ,       �        ���������                                4       �	        ���������	                                4       �	        ,   �����	        ���������	            �		�	�	�	�	4	 	�	�	                        4       4	��@ ,   ����4	 � ��������4	  � ios_base::_M_grow_words is not valid    ios_base::_M_grow_words allocation failed St8ios_base   �			        		�"0#                                            J   �    @                     �   @                      -+xX0123456789abcdef0123456789ABCDEF -+xX0123456789abcdefABCDEF -0123456789 GMT HST AKST PST MST CST EST AST NST CET IST EET JST     locale::_S_normalize_category category not found    locale::_Impl::_M_replace_facet p) )`)P)@)0)NSt6locale5facetE   �	�
	        �
	p$�$C   ?                              St15basic_streambufIcSt11char_traitsIcEE    �	 	                ,	202`1p1�1�1�1�1@3�1 3�1`2 2basic_ios::clear                St9basic_iosIcSt11char_traitsIcEE   	�			    �	�:�:St7codecvtIcc9mbstate_tE    	�	��                            �	�C0D@C`CpC�C�C�C�Cbasic_filebuf::underflow codecvt::max_length() is not valid basic_filebuf::underflow incomplete character in file   basic_filebuf::underflow invalid byte sequence in file  basic_filebuf::underflow error reading the file basic_filebuf::xsgetn error reading the file    basic_filebuf::_M_convert_to_external conversion error                  St13basic_filebufIcSt11char_traitsIcEE  	�	,	            St14basic_ifstreamIcSt11char_traitsIcEE 	�	�	            St14basic_ofstreamIcSt11char_traitsIcEE 	 	�            St13basic_fstreamIcSt11char_traitsIcEE  	`	�	                                                �	�a�w�] H�Z�\ I�H P�K 30I�J�Xh       �	        ���������	        L		 	`	        h       	Py�z��������	�y@{                        d       �        ���������        �	�	�	�	        d       H	�xPz��������H	@y�z                        d       �        ���������                                l       �	        ���������	                                l       �	        d   �����	        ���������	            	�	L	`		 	�	�	4	 	                        l       �	P{�{d   �����	�{@|���������	�{P|basic_string::at: __n (which is %zu) >= this->size() (which is %zu) basic_string::_S_construct null not valid basic_string::copy basic_string::compare basic_string::_S_create basic_string::_M_replace_aux basic_string::insert basic_string::replace basic_string::assign basic_string::append basic_string::resize basic_string::basic_string basic_string::substr   ���?����std::future_error regex_error St11regex_error   	�	$	    �	 �0��std::bad_cast St8bad_cast   	
	�	        	����p�    N10__cxxabiv121__vmi_class_type_infoE   	@	d	                h	��ж������`�`�� �std::exception std::bad_exception St9exception  �	�	St13bad_exception   	�	�	                            N10__cxxabiv115__forced_unwindE �	 	                        N10__cxxabiv119__foreign_exceptionE �	`	        �	 �`�@�        �	0�p�P�        @	        ��        �	        ��St9type_info    �	�	                                �	�� ��������N10__cxxabiv117__class_type_infoE   	@	�	                    d	����������`� ����std::bad_alloc St9bad_alloc 	�	�	        �	������std::bad_typeid St10bad_typeid  	�	�	    	0�@� �                    N9__gnu_cxx20recursive_init_errorE  	@	�	    d	p���@�pure virtual method called
 deleted virtual method called
  N10__cxxabiv120__si_class_type_infoE    	�	d	                �	����������`����� �terminate called recursively
 '
   what():      terminate called after throwing an instance of '    terminate called without an active exception
 std::bad_array_length St16bad_array_length    	�	�	    �	������l	\	T	D	0	(	    �E    �E�E�E�E    �E�E�E    �E    �E�E�E    �E�E    NSt8ios_base7failureE   	x	�	        �	������Sd          �	�	      �	   �         �        ���������                                       �	        ���������	        �	,	@	�	 	�	�	                                   �	�� �   �����	��0����������	��@�true false Si   �	�	       �	���    	 	                       �	�� ����������	��@�ab a+ rb a+b wb r+ r+b w+ w+b                                                           �7	            (	        �	+	        .	1	        y8	�7	        5	(	        8	+	        ;	1	                                                                        y8	            5	            ?	            B	St11logic_error 	p	�	St12domain_error    	�	�	St16invalid_argument    	�	�	St12length_error    	�	�	St12out_of_range    	�	�	St13runtime_error   		�	St11range_error 	0	$	St14overflow_error  	L	$	St15underflow_error 	l	$	        �	���        �	� �        �	0@�        �	p��        	���        $	 �        @	`p�        `	���        �	���%Lf LC_CTYPE LC_NUMERIC LC_TIME LC_COLLATE LC_MONETARY LC_MESSAGES  locale::facet::_S_create_c_locale name not valid    h	q	|	�	�	�	�	������������������������������      ���������      AM PM Sunday Monday Tuesday Wednesday Thursday Friday Saturday Sun Mon Tue Wed Thu Fri Sat January February March April May June July August September October November December Jan Feb Mar Apr Jun Jul Aug Sep Oct Nov Dec bad_function_call St17bad_function_call    		�	        8	�!�!p!not enough space for format expansion (Please submit full bug report at http://gcc.gnu.org/bugs.html):
     future Broken promise Future already retrieved Promise already satisfied No associated state Unknown error              *N12_GLOBAL__N_121future_error_categoryE    	@ 	�!	St12future_error    	x 	�	            l 	�#�#�#�%`'�(�'        � 	$ $P$generic system                      *N12_GLOBAL__N_122generic_error_categoryE                       *N12_GLOBAL__N_121system_error_categoryE    	@!	�!		 !	�!	St14error_category  �	�!	St12system_error    	�!	$	    x!	�'�'@' (`'�(�'                                l!	�'�'P'�'`'�(�'                                �!	        ����`'�(�'        �!	P(`(� std::bad_array_new_length St20bad_array_new_length 	�"	�	        �"	�)�)�)                                            `*P*P*P*P*`*`*`*`***P*************`*********P******`***T*P*`*P***T*`*`***P*P*P*P*P**P*P**P*`*`****`*`*`****P*P*G.k.k.k.�.G.G.@.@.k.k.k.k.k.k.k.k.k.k.k.k.k.k.k.G.k.k.k.k.k.k.k.k.k.k.`.`.k.k.G.k.k.k.k.k.k.k.k.k.G.@.k.k.k.k.k.k.k.k.k.k.k.k.G.G.k.P.P.P.P.G.k.k.k.k.k.�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�2�GCGCGH�EcE�D�D�DD^D#DD�C�C�C~CJ�I�I�IK�J�FIFMJMJMJ@J@J@J@J@J@J@JII@J@J�HiC'C�A�A?�A>>�>=�=�<�<D<�?�?�@V?V?|5|5e?!<�;�:#:�9#9�8$Ku8s;T8X77�6�V�V�V�V�V�]]]]]]]]]]]]]]]]]]]]]]�]@^�^�]@^�^@_�_�\@`�`�`�` a]]]]�a]0]P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�`�P���0�P�� �P�P�P�P�P�`�P����P��@�0���P�P�P�P�P�P�P�P�P�P�P�����������P�����P�P�P���������U�P�P�P�P�P�P�P�P�P�P�P�P�P�d�P�P�P�P�P�P�P�P�P�P�P�P�?�P�P��)���P���~�P�P�P�P���P���P�P�n�d�P�b����� �� �:���������P�@�@�P�P�P�P�����P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�P�����z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�p�z���z�@�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�z�`���z�z�h�z�F����z�z�z�z�z�z�z�z�����z�z�X�z�z�z�z�z�z�z�z�z�z�z��z�z�z�z���z�z�z�z�z�z�z�z�z�z�z�z�z��t   (7	   (7	           a   ,7	   ,7	   17		   b   ;7	   ;7	   @7	   s   M7	   �9	F   @7	   i   Y7	   0:	1   f7	   o   t7	   d:	1   �7	   d   �7	   �:	2   �7	                                                               �7	�7	      �7	p8	      �7	�6	      "6	�6	      �	�6	      �	�7	      �7	�7	      �7	�7	
      (6	�7	      �7	�7	      �7	�7	      �7	�7	      �7	�7		      �7	�7	      8	8	      8	8	      8	8	      7	Z6	      8	8	      8	8	      !8	$8	      &8	)8	      ,8	�8	      %6	�4	      /8	�8	      +6	l8	      28	58	      9	68	      7	98	      E8	H8	      K8	I8	      N8	Q8	      T8	W8	      Z8	d8	      ]8	8	      `8	c8	      f8	i8	      �	o8	      V7	d8	      B9	r8	      t8	w8	      {8	~8	      �8	�8	      0 	�8	      �8	�8	      �8	�8	      �8	�8	      �8	�8	      �8	�8	      7	�8	      .6	�8	      �8	�8	      �8	�8	      �8	�8	      �8	�8	      �8	�8	      �8	�8	      �7	�8	      �8	�8	      �	�8	       �8	�8	                                                      ,9	   ,9	       �8	    9	      39	   9	       9	   9	      9	   9	      9	   9	      9	
   9	
      *9	   *9	       A9	   A9	      89	   E9	                          W9	   W9	      N9	   N9	      e9	   e9	       \9	   \9	                                                                   w9	   w9	       n9	   n9	                           }9	   }9	   	   �9	   39	       �9		   W9	      �9	   �9	      X6	   X6	       �9		   �9		       �9		   �9		       �9	
   �9	
       �9	   �9	      �9	   �9	       �9	   �9	       �9	   �9	       _GLOBAL_ (anonymous namespace) %ld [abi: {default arg# }:: JArray VTT for  construction vtable for  -in- typeinfo for  typeinfo name for  typeinfo fn for  non-virtual thunk to  covariant return thunk to  java Class for  guard variable for  TLS init function for  TLS wrapper function for  reference temporary # hidden alias for  non-transaction clone for  _Sat  _Accum _Fract ,  operator operator  ad gs cl ix qu  :  new  ull java resource  decltype ( ... this {parm# global constructors keyed to  global destructors keyed to  {lambda( )# {unnamed type#  [clone  >(  restrict  volatile  const && complex  imaginary  ::*  __vector( dt pt auto li string literal std std::allocator std::basic_string std::string std::istream basic_istream std::ostream basic_ostream std::iostream basic_iostream aN &= aS aa alignof  az cc const_cast () cm , co ~ dV /= da delete[]  dc dynamic_cast de dl delete  ds .* dv / eO ^= eo ^ eq == ge gt lS <<= operator""  ls << lt mI -= mL *= mi ml mm -- na new[] != ! nw new oR |= oo || pL += pl pm ->* pp ++ ps -> ? rM %= rS >>= rc reinterpret_cast rm % rs >> sc static_cast sizeof  sz throw tw throw  bool boolean byte long double float __float128 unsigned char unsigned int unsigned unsigned long unsigned __int128 unsigned short void wchar_t unsigned long long decimal32 decimal64 decimal128 half char16_t char32_t decltype(nullptr)    std::basic_string<char, std::char_traits<char>, std::allocator<char> >  std::basic_istream<char, std::char_traits<char> >   std::basic_ostream<char, std::char_traits<char> >   std::basic_iostream<char, std::char_traits<char> >  d�������&���E���d����������F�������Ư��?���r����������E���{���Ʊ��6��������������������}���}���}���}���}���}���}���}���}���}���}���}���}���}���}���}���}���}���}���}���}���}���d�������f���ٴ��)��� ���ٴ�����}���}���}���}���X���k���ٴ��������b���Y������?���D���D���D���D��������������?����������\����������D���D���D���D���i���������������������������������Խ��Ľ������������������4���4�������������������������������d����������$���$���$���$���$���������$���$������$���$���$���$�������$���$���$���$���$���$��������������������������������������������������������������������������������������������������������������������������������������D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���D���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���4���ľ������$������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������������4������� �����������F�������������������������������F���S���\���j���s���������������������������(���1���:�������C�����������������������������������������d���T����������T���������������������������T�������                                            ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                            failed to parse command line arguments C                                            ��������                                                                                                                                                                                                                                                                            max system bytes = %10lu
 system bytes     = %10lu
 in use bytes     = %10lu
                                               ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                            '"sscanf"' is not implemented                                               ��������                                                                                                                                                                                                                                                                            r w                                                 ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                            '"strtod"' is not implemented                                               ��������                                                                                                                                                                                                                                                                          �'"strtof"' is not implemented                                               ��������                                                                                                                                                                                                                                                                          �                                            ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                            '"strcoll"' is not implemented                                              ��������                                                                                                                                                                                                                                                                            ERROR(TODO)                                                 ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                            warning: fstat(%i, %x) not implemented                                              ��������                                                                                                                                                                                                                                                                            warning: strftime("%s") is not implemented                                          ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                    0123456789abcdef 0123456789ABCDEF 012345678 0123456789   - + 0 x X .    =�Z�Z�G�Z�Z�Z�Z�Z�Z�Z�3�Z�)�Z�Z�Q�^�y�y�y�^�^�^�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y�y� �y�y�y�y�y�y�y�y�^�y�&� �^�^�^�y� �y�y�y�y�[� � �y�y���y� �y�y� �-�D�^�v��������� �:�W�t���������                                                ��������                                                                                                                                                                                                                                                                                           �>@            $@      �C                                            ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                                                                        ��������                                                                                                                                                                                                                                                                               zR |�        ����
    A�BF�     <   ����    A�BI�         zPLR |  � �  <   $   *����  D Gu Duxu|W.� A�A�C   ,   d   p���E  >A�BD�.*��      �   ����$   A�B �     ����@    A�B|�     ,  �����    A�B}�    L  
���L    A�BH�    l  6���A    A�B}�     �  W���    A�BV�     �  ^���
    A�BF�  (   t  H����   iA�BD�_.���     �  ѓ���    A�B��      H���A    A�B}�     8  i���    A�BV�     X  c���
    A�BF�     x  M���A    A�B}�     �  n���    A�BV�     �  h���
    A�BF�  (   �  R���3  {A�BG�}.���      Y���A    A�B}�     $  z���    A�BV�     D  t���
    A�BF�      d  ^���0    A�BD�h��     �  j���     A�B\�     �  j���c    A�B_�    �  ����
    A�BF�  (   �  ����  �A�BD��.Z��      x���    A�BY�     4  v���    A�BZ�     T  t���    A�B[�     t  t���     A�B\�     �  t���    A�BX�     �  p���    A�BS�     �  t���       (   �  p���@    A�A�C�x�A�A�D     ����K    A�A�C�G,I0F P$G(A,A0F MA�A�A� P   \  ����   A�A�C�A�E@M
C�A�A�A�B�C�A�A�A� (   �  H����    A�C j,M0LA�H � P   �  ����s    A�A�C�A�E0Y
A�A�A�A�ACC�A�A�A�  @   0  ؗ��p    C\A HC
EE
KSA HC
ACA HCP   t  ���   A�A�C�A�G0K<A@H0h<C@L0�
A�A�A�A�I   �   p  �����  �A�A�F�A�Cpb
A�A�A�A�NetGxB|G�HtAxB|G�F|AxA|G�HpH
A�A�A�A�F]|G�LprxI|G�Hpi|E�QpL|I�QpL|K�Jp�
|G�O|A�Tph|A�  0   H  ����   �A�BF���_.k. Q.L. h. $   |  ����*   �A�BF.I
�A8   �  ����P    A�C_A EG
A�OC
A�ACC    8  ����c    A�C~O      X  ���V    A�CrA P  (   |  ,���E    A�CK
A XMC H    �  P���          �  L���          �  X���           �  T���+    A�CU LA�    	  `���          	  \���%       4   �  x����   �A�BF���S.L
�A�A�A�A     h	  О��          |	  ܞ��           �	  ؞��    A�CL GC�     �	  Ԟ��    A�CL GC� @   �	  О��V    A�A�CTDA FZ
A�A�PCA�A� 4   �	  ����   A�BD�V.Q
��B`
��A`. <   �	  �����   DA�BE��f
�A�A�PU. ^
�A�A�C`. 8   <
  4����   |A�BF���V
�A�A�A�Nd. M.    8   x
  �����   �A�BF���\
�A�A�A�HT. M.         ����%       4   �
  ȡ���   �A�BF���R.L
�A�A�A�A  <   X   ���e    A�A�ChA HT
A�A�DNA�A�H   �  P���a    A�A�CgC FH
A�A�AFLA HCA�A�D   �  t���T  A�BC���u.\
�A�A�A�Fq
�A�A�A�A|.  D   �  ����i  HA�BC���l
�A�A�A�Ka
�A�A�A�LL.T. D     ����B  �A�BC���o.[
�A�A�A�Ma
�A�A�A�A`.     �  ����       L   �  ����s    A�A�C^AA LA�A�M��CA JSBA E        ���    CBD H      @  ���       P   T  ���z    A�A�A�\
�A�A�O\
�A�A�BCA JMBA E    �  ���          �  ���          �  (���G    A�u
�J      �  X���            d���       P   �  p���   �A�BI����
�A�A�A�HR.�
�A�A�A�L�. O.@.       l  ���    C$J(E,D0H   �  ���    C$J(E,D0H   �  ���    C$J(E,D0HT   �  ���R    A�A�COA HAAA HE
A�A�AELA HEA�A�T   $  $���R    A�A�COA HAAA HE
A�A�AELA HEA�A�T   |  ,���R    A�A�COA HAAA HE
A�A�AELA HEA�A�H   |  4���  A�BI���X. ^.
�A�A�A�La
�A�A�A�LB.       ����          4  ����@          H   ���       H     ���  TA�BI���X. ^.
�A�A�A�La
�A�A�A�LB.    �  ���          �  ܭ��          �  ح��       H   �  ԭ��  �A�BF���p. ^.
�A�A�A�Ga
�A�A�A�LB.    0  ����       H   �  ����  �A�BF���g. ^.
�A�A�A�Pa
�A�A�A�LB.    �  x���       H   L  t���  ,A�BF���g. ^.
�A�A�A�Pa
�A�A�A�LB.    �  H���       H   �  D���  tA�BI���^. ^.
�A�A�A�Fa
�A�A�A�LB.    P  ���          d  ���    CK H  H   (  ���  �A�BI���^.0^.
�A�A�A�Fa
�A�A�A�LB.    �  ̶��       H   �  ȶ��  A�BI���X. ^.
�A�A�A�La
�A�A�A�LB.    ,  ����          @  ����           T  ����$    A�CN LA�     x  ����    A�CG KA� ,   �  ����     A�CG FACA HA� ,   �  ����?    A�CPCA HJ
A�E    �  ����       @     ����j    A�A�HoAAC HGC MFC�A�       T  ĸ��    CGDBD H D   x  ����M    A�A�CKDBA HO
A�A�PJA�A�      �  ȸ��I    C[
RCC M t   �  �����    A�A�C`OAC HG
C�A�ECC HK
C�A�CCDB A$A(A,A0B,CEA�A�   \  ���    CIAD HP   |  ���s    A�A�C^ADA HA�A�M��CA JSBA E       �  8���Z    A�Cx \A�    �  t���       H   �  p���  LA�BI���h
�A�A�A�IJ
�A�A�A�C�.�.   H   �  4����  �A�BF���0
�A�A�A�Di.f
�A�A�A�A�.   <   H  ����  �A�BI���H.�
�A�A�A�F�.    8   �  ����X  8A�BI���K
�A�A�A�AO.a.  8   �  ����  �A�BI���~
�A�A�A�CO.H.      X  ����          l  ����          �  ����          �  ����          �  ����          �  ����          �  ����          �  ����          �  ����            ����             ����          4  ����          H  ����          \  ����          p  ����          �  ����          �  ����          �  ����          �  ����          �  ����!    A�_�     �  ����            ����            ����          ,  ����          @  ����          T  ����          h  ����          |  ����          �  ����       (   �  ����&    A�C$I(J,A0HC�   (   �  ����&    A�C$I(J,A0HC�   (   �  ����&    A�C$I(J,A0HC�   (   (  ����&    A�C$I(J,A0HC�   (   T  ����&    A�C$I(J,A0HC�   (   �  ����&    A�C$I(J,A0HC�   (   �  ����&    A�C$I(J,A0HC�   (   �  ����&    A�C$I(J,A0HC�   (     ����&    A�C$I(J,A0HC�   (   0  ����&    A�C$I(J,A0HC�   (   \  ����&    A�C$I(J,A0HC�   @   �  ����m    A�CZA HJA HJA HJA HGA�@   �  ����m    A�CZA HJA HJA HJA HGA�8     ���Z    A�CZA HJA HJA HGA�     L  ,���    A�CE LA�     p  (���    A�CE LA�     �  $���!    A�CK LA�     �  0���!    A�CK LA�     �  <���!    A�CK LA�        H���!    A�CK LA�     $  T���    A�CE LA�     H  P���!    A�CK LA�     l  \���!    A�CK LA�     �  h���!    A�CK LA�     �  t���    A�CE LA�     �  p���!    A�CK LA�     �  |���!    A�CK LA�        ����!    A�CK LA�     D  ����!    A�CK LA� (   h  ����"    A�CMAD HC�   0   <  ����>   �A�BB��P.O
�A�A�E       �  ����    A�CE LA�    �  ����              ����!    A�CK LA� 0   �  ����>   �A�BB��P.O
�A�A�E   0      ����m   �A�BB��r.\
�A�A�E       �  ����    A�CE LA�    �  ����           �  ����!    A�CK LA� 4   �   ���2    A�CP
A�KCAA HCA�  D   �  ���'  A�BI���e.{
�A�A�A�AB
�A�A�A�K   H   h   ����@    A�A�GA JM
C�A�KCAA ECA�A�   0   \   ����>   A�BB��P.O
�A�A�E   0   �   ����F   *A�BB��P.W
�A�A�E   0   �   ���F   :A�BB��P.W
�A�A�E   H   �   (����  LA�BI���T.
�A�A�A�CN
�A�A�A�CQ.    �   �!  �����    A�A�F�CBB YKADD HE
�A�A�ECA SCAA FAEB LADD FAAB RC�A�A� l   ,"  �����    A�A�A�A�C n$C(A,A0HC�A�A�A�H ����C,A0J ]A�A�A�A�  �   �"  ����(   A�A�A�A�C0_
A�A�A�A�FL<A@H0V
C�A�A�A�Oc<A@H0i<A@H0i<A@H0S<A@H0W<A@H0g<A@H0g<A@H0W<A@H0W<A@H0 0   �"  l���L   xA�DB��c.L
�A�A�A   0   (#  ����K   �A�DB��b.L
�A�A�A   0   \#  ����N   �A�DB��e.L
�A�A�A      �#  ����"          �#  ����"       D   $  ����S    A�C X$E(F,A0H E
A�JC(A,A0B,C EA�D   X$  ���S    A�C X$E(F,A0H E
A�JC(A,A0B,C EA�D   �$  (���S    A�C X$E(F,A0H E
A�JC(A,A0B,C EA�D   �$  @���S    A�C X$E(F,A0H E
A�JC(A,A0B,C EA�   0%  X���"       (   D%  t���H    C `
MC(A,A0F,C G(   p%  ����H    C `
MC(A,A0F,C G0   D%  ����L   �A�DB��c.L
�A�A�A   0   x%  ����K   �A�DB��b.L
�A�A�A   0   �%  ����N   �A�DB��e.L
�A�A�A      8&  ���"          L&  ,���"       D   `&  H���S    A�C X$E(F,A0H E
A�JC(A,A0B,C EA�D   �&  `���S    A�C X$E(F,A0H E
A�JC(A,A0B,C EA�D   �&  x���S    A�C X$E(F,A0H E
A�JC(A,A0B,C EA�D   8'  ����S    A�C X$E(F,A0H E
A�JC(A,A0B,C EA�   �'  ����"       (   �'  ����H    C `
MC(A,A0F,C G(   �'  ����H    C `
MC(A,A0F,C G   �'  ����           (  �����       @   �'  ����   �A�DF���`.t
�A�A�A�Nn
�A�A�A�A @    (  �����   �A�DF���`.t
�A�A�A�Nn
�A�A�A�A    �(  ���       @   �(  (���>    A�CND D$F(D,D0D4D8A<A@C<CC�   @   �(  $���>    A�CND D$F(D,D0D4D8A<A@C<CC�      8)   ���       @   L)  ,���@    A�CND D$F(D,F0D4D8A<A@C<CC�   8   �)  (���8    A�CNFDF D$D(A,A0C,CC� 0   t)  ,���J   �A�DB��a.L
�A�A�A   0   �)  H���I   �A�DB��`.L
�A�A�A   0   �)  d���K   A�DB��b.L
�A�A�A      h*  ����"          |*  ����"       D   �*  ����S    A�C X$E(F,A0H E
A�JC(A,A0B,C EA�D   �*  ����S    A�C X$E(F,A0H E
A�JC(A,A0B,C EA�D    +  ����S    A�C X$E(F,A0H E
A�JC(A,A0B,C EA�   h+   ���S       @   $+  L����   A�DF���^.t
�A�A�A�Pk
�A�A�A�A    �+  ����       <   �+  ����8    A�CN D$D(D,D0D4D8A<A@C<CC�  <   ,  ����8    A�CN D$D(D,D0D4D8A<A@C<CC�  <   T,  ����8    A�CN D$D(D,D0D4D8A<A@C<CC�  <   �,  ����8    A�CN D$D(D,D0D4D8A<A@C<CC�  <   �,  ����8    A�CN D$D(D,D0D4D8A<A@C<CC�     -  ����       4   (-  ����4    A�CPFD D$D(A,A0C,CC�8   `-  ����6    A�CNDFD D$D(A,A0C,CC� <   �-  ����:    A�CN D$D(F,D0D4D8A<A@C<CC�  4   �-  ����2    A�CNFD D$D(A,A0C,CC�0   �-  ���R   ,A�DB��i.L
�A�A�A   0   �-  0���Q   8A�DB��h.L
�A�A�A   8   $.  \����   DA�DF���@.L
�A�A�A�Fq.      �.   ���          �.  ���          �.  ���          �.  $���          /   ���          /  ,���G          0/  h���G          D/  �����          X/   ����          l/  �����         �/  8���       <   �/  D���>    A�CP F$D(F,D0D4D8A<A@C<CC�     �/  D���          �/  P���          �/  \���       <   0  X���8    A�CN D$D(D,D0D4D8A<A@C<CC�  <   P0  X���8    A�CN D$D(D,D0D4D8A<A@C<CC�  <   �0  X���8    A�CN D$D(D,D0D4D8A<A@C<CC�  <   �0  X���8    A�CN D$D(D,D0D4D8A<A@C<CC�  <   1  X���8    A�CN D$D(D,D0D4D8A<A@C<CC�     P1  X���       4   1  d���>   dA�A�Ea
A�A�AEA   4   D1  l���>   pA�A�Ea
A�A�AEA      �1  t���          �1  p���       4   �1  l���,    A�CND D$D(A,A0C,CC�      42  d���          H2  `���          \2  \���       @   2  X����   |A�BC���F
�A�A�A�AG.Z
�A�A�A�A@   \2  �����   �A�BC���F
�A�A�A�AG.Z
�A�A�A�A4   �2  ����>   �A�A�Ea
A�A�AEA       03  ����.    A�E[ KA�    T3  ���       ,   h3   ���$    A�CNDAA CCC�    �3   ���       @   T3  �����   �A�DF���H
�A�A�A�JG.Z
�A�A�A�A,   �3  h���L    CE LSEEA HG
A �    4  �����   A�A�A�A�CLbPH@�LKPATDXD\D`DdDhDlEpCld@m
C�A�A�A�M�DBHALAPE@[DBHALAPE@`DBHALAPI@_HGLAPF@ x   �4  ����   A�A�A�A�HL`PL@�
A�A�A�A�G3LCPF@^DBHALDPE@MLCPF@{LGPJ@kLCPF@  �   @5  H���X   A�A�A�A�CLTPT@EDAHBLEPBTEXD\D`AdAhDlApElK@T
A�A�A�A�FyLAPF@CLCPF@  ,   �5  $���L    CE LSEEA HG
A ,   �5  D���L    CE LSEEA HG
A ,   $6  d���L    CE LSEEA HG
A H   �5  ����M  �A�BF���u.�
�A�A�A�Es
�A�A�A�J�.  ,   �6  ����L    CE LSEEA HG
A ,   �6  ����L    CE LSEEA HG
A ,    7  ����L    CE LSEEA HG
A H   �6  �����  HA�BF����.
�A�A�A�Ho
�A�A�A�Ng.  ,   |7  ,���L    CE LSEEA HG
A H   T7  L����  �A�BF����.
�A�A�A�Ho
�A�A�A�Ng.  ,   �7  ����L    CE LSEEA HG
A ,   (8  ����L    CE LSEEA HG
A ,   X8  ����L    CE LSEEA HG
A ,   �8  �����   A�BI���
�A�A�A�J,   �8  `���L    CE LSEEA HG
A ,   �8  ����L    CE LSEEA HG
A ,   9  ����L    CE LSEEA HG
A 4   H9  ����I    A�CE NUEEA HHA�   4   �9  ����I    A�CE NUEEA HHA�   4   �9  ����I    A�CE NUEEA HHA�   4   �9  ���I    A�CE NUEEA HHA�   4   (:   ���I    A�CE NUEEA HHA�   4   `:  8���I    A�CE NUEEA HHA�   4   �:  P���I    A�CE NUEEA HHA�   4   �:  h���I    A�CE NUEEA HHA�   4   ;  ����I    A�CE NUEEA HHA�   4   @;  ����I    A�CE NUEEA HHA�   4   x;  ����I    A�CE NUEEA HHA�   4   �;  ����I    A�CE NUEEA HHA�   4   �;  ����I    A�CE NUEEA HHA�   <    <  �����   A�A�C�A�C x
A�A�A�A�K�   `<  h����    A�A�A�A�C _(F,A0F4A8A<A@J$K(A,A0J G
A�A�A�A�NE(F,A0D4A8A<A@H GA�A�A�A�   8   �<  x���5    A�A�CQA D$D(F,A0LA�A� P   �<  |���  �A�BF����.F. s.Z. [.X. _.^
�A�A�A�Jv. S.P   (=  H��  �A�BF����.F. s.Z. [.X. _.^
�A�A�A�Jv. S.D   |=  ���  H A�BC���b.Y. _. S.y. f
�A�A�A�Kd.   d   >  ���w    A�CZGAA D$D(A,A0E,CE
A�QCGAA D$D(A,A0E,CEA�  �   �>  ���4   A�A�A�A�C0}4A8F<A@^A�A�A�A�R0����C<D@H0d4A8A<C@YA�A�A�A�K0����c<A@P0�8B<A@I08    ?  h��/    A�A�CJA D$D(F,D0JA�A� 4   \?  \���    A�A�A�A�
�A�A�A�A8   <?  ���  ` A�BF���K
�A�A�A�I�.�. H   x?  ����  � A�BF���m
�A�A�A�G�
�A�A�A�P�.�.   4   @  L��1    A�CHFD D$D(D,A0E,CC�p   T@  T��r    A�A�CaDAA D$D(A,A0E,CE
A�A�KCDAA D$D(A,A0B,CEA�A� 8   p@  `���  � A�BF���
�A�A�A�H�.�. 4   A  ���1    A�CHFD D$D(D,A0E,CC�T   <A  ���p    A�A�A�A�C0e4D8F<A@ADAHDLAPELfA�A�A�A�  p   �A  ���r    A�A�CaDAA D$D(A,A0E,CE
A�A�KCDAA D$D(A,A0B,CEA�A� X   B  ���   A�A�A�A�C0k4B8L<A@M0D4B8A<A@J0S
C�A�A�A�A8   B  ���(  � A�BF���f
�A�A�A�N�.�. 8   �B  ���5    A�CHDFD D$D(D,A0E,CC� �   �B  ���o    A�A�A�A�C g$A(A,A0D4D8A<A@E<C E
A�A�A�A�DA$A(A,A0D4D8A<A@B<C EA�A�A�A�   8   C  ����  !A�BF���+
�A�A�A�I�.�. 8   �C  !��5    A�CHDFD D$D(D,A0E,CC� �   �C  !��o    A�A�A�A�C g$A(A,A0D4D8A<A@E<C E
A�A�A�A�DA$A(A,A0D4D8A<A@B<C EA�A�A�A�   H   D  � ��(  L!A�BF���d
�A�A�A�PE.�
�A�A�A�AP. V.  H   hD  �!��(  t!A�BF���d
�A�A�A�PE.�
�A�A�A�AP. V.  H   �D  �"���   �!A�BF���d
�A�A�A�PE.o
�A�A�A�AP. V.  ,   XE  p#���   A�BC����
�A�A�A�D<   �E   &��7    A�CH D$B(F,D0D4D8D<A@E<CC�  ,   �E   &���   A�BC����
�A�A�A�J@   �E  �(��;    A�CHD D$B(F,D0D4D8D<A@E<CC�   <   <F  �(��c    A�CU
A�FQ
A�NCC FN
A�AX   |F  �(���    A�A�C t
A�A�Ex
A�A�FC,C0F ],A0F ]
A�A�A  ,   �F  �)��   A�BF���a
�A�A�A�C ,   G  p,���   A�BC����
�A�A�A�I�   8G  @0��   A�A�A�A�C|V��tExG|B�E�E�G�G�G�G�G�A�E�gpK
A�C�A�A�Fy|A�FpC|C�Fp   �   �G  �1���   A�A�A�A�F�Y�G�E�G�B�E�E�G�G�G�G�G�A�E�g�N
A�C�A�A�Jy�A�F�C�C�F� �  `H  4��=   A�A�A�A�C|K�R|G�Jp�|C�Fp~
A�A�A�A�RY|A�FpGtBxA|A�EpfxC|N�E�G�G�G�G�G�G�E�E�[pH|H�Kpm|H�Kpd|A�ZpPtGxB|B�B�E�G�G�G�G�G�E�E�Ypv|H�HtDxB|A�Hp]|A�SpE
tGxB|B�B�A�JEtGxB|B�B�K�J�G�G�G�G�E�E�SpF
xC|G�tExG|B�E�K�G�G�G�G�G�E�E�LpC
tExG|B�E�ZC|H�HtDxB|A�HpKtExG|B�E�E�G�G�G�G�G�E�E�YxH|H�Hpc|H�LpW|H�LpYtGxB|B�B�E�G�G�G�G�G�E�E�YpAtGxB|B�B�E�G�G�A�A�G�E�E�YpS
xC|GE
tExE|A�F|AxA|HE
tGxB|B�B�G�GE
tExE|A�F|AxA|HE
tGxB|B�B�K�SE
tGxB|B�B�K�SE
tGxB|B�B�K�SE
tExE|A�F|AxA|HEtGxB|E�B�E�G�G�G�G�G�E�E�Yp)|A�FpztBxA|A�EpN
tGxB|B�B�K�EUtExA|A�EpH|C�FpHtExA|A�EpGtExA|A�Epx   @L  h=��   A�A�A�A�C<T@O8C<D@DDAHDLDPATAXD\A`E\K0w
A�A�A�A�Pj<C@F0u<A@F0  x   �L  >��   A�A�A�A�C<T@O8C<D@DDAHDLDPATAXD\A`E\K0w
A�A�A�A�Pj<C@F0u<A@F0  L   �L  �>���  �!A�BF���T.�
�A�A�A�Ep. t.�
�A�A�A�CL   0M  L���  �!A�BF���T.�
�A�A�A�Ep. t.�
�A�A�A�C8   �M  pY���   �!A�BI���m.0N. z
�A�A�A�LW.0 8   �M  $Z���  "A�BF���.0B
�A�A�A�Cy.   D   �M  �[���
  "A�BC����.�
�A�A�A�JE	
�A�A�A�C <   @N  Pf��k  A"A�BC���S.a.0T. k
�A�A�A�Dh. <   �N  �g��k  P"A�BC���S.a.0T. k
�A�A�A�Dh. <   �N  �h��k  _"A�BC���S.a.0T. k
�A�A�A�Dh. D    O  �i���  n"A�BF���/
�A�A�A�EL.
�A�A�A�C <   �O  hr��7    A�CH D$D(D,D0D4D8D<A@E<CC�  p   �O  hr��|    A�C\D D$A(D,D0D4D8A<A@E<CE
A�GCD D$A(D,D0D4D8A<A@B<CEA�  �   TP  tr��d   A�A�A�A�C@]LEPDTAXD\D`DdDhDlApElW@PHRLEPH@eHILEPM@LCPF@GLCPF@K
A�A�A�A�MiLAPF@KLCPF@ D   �P  @v���  �"A�BF���&
�A�A�A�NL.
�A�A�A�C <   @Q  �~��7    A�CH D$D(D,D0D4D8D<A@E<CC�  p   �Q  �~��|    A�C\D D$A(D,D0D4D8A<A@E<CE
A�GCD D$A(D,D0D4D8A<A@B<CEA�  D   �Q  �~���  �"A�BF���&
�A�A�A�NL.�
�A�A�A�C <   <R  \���7    A�CH D$D(D,D0D4D8D<A@E<CC�  p   |R  \���|    A�C\D D$A(D,D0D4D8A<A@E<CE
A�GCD D$A(D,D0D4D8A<A@B<CEA�  D   �R  h����  �"A�BF���&
�A�A�A�NL.�
�A�A�A�C <   8S  ����7    A�CH D$D(D,D0D4D8D<A@E<CC�  P   xS  ����l    A�A�A�C0O<S@DDAHDLDPDTDXD\A`E\_A�A�A� p   �S  ����|    A�C\D D$A(D,D0D4D8A<A@E<CE
A�GCD D$A(D,D0D4D8A<A@B<CEA�  D   �S  ����	  �"A�BF����
�A�A�A�G\.d
�A�A�A�C <   �T  ����7    A�CH D$D(D,D0D4D8D<A@E<CC�  p   �T  ����|    A�C\D D$A(D,D0D4D8A<A@E<CE
A�GCD D$A(D,D0D4D8A<A@B<CEA�  D   �T  ̙���	  �"A�BC���W
�A�A�A�PL.�
�A�A�A�C <   �U  4���7    A�CH D$D(D,D0D4D8D<A@E<CC�  p   �U  4���|    A�C\D D$A(D,D0D4D8A<A@E<CE
A�GCD D$A(D,D0D4D8A<A@B<CEA�     8V  5���          LV  ,���          `V  (���          tV  $���          �V   ���          �V  ���          �V  ���       0   lV  ���W   �"A�BB��P.h
�A�A�E       �V  @���    A�CE LA� (   W  <���"    A�CMAD HC�   �   HW  @���    A�A�C�A�F�k�L�A�A�H�Q
A�A�A�A�A\
A�A�A�A�AC�A�F�H�A�A�E�I�E�B�E�A�A�J�  d   �W  �����    A�A�C�A�F�^�I�A�A�H�N
A�A�A�A�AA�L�A�A�E�,   �W  ����  #A�BD��.�
��A   �X  ����%       ,   @X  ����_   4#a�BH.a
�AM�   ,   pX  ���F  H#A�BD��.�
��B  0   �X  ���m   \#A�BB��M.c
�A�A�E       ,Y  L���    A�CE LA� 8   PY  H���l    A�C V
A�Ec$B(A,A0K C
A�J    �Y  |���    A�CE NA� @   XY  x����   l#A�BF���u
�A�A�A�OM.u
�A�A�A�A @   �Y  ����   ~#A�BF���].X
�A�A�A�OB
�A�A�A�A   8Z  P���
          LZ  L���
       �   `Z  H���   A�A�A�A�C y$D(A,A0F L,C0F R
C�A�A�A�Gs(G,A0F O
C�A�A�A�JC,C0F W,E0F      �Z  ܪ��6           [  ���F       <   [  D���W    A�A�A�u
�A�A�FI
�A�A�E  ,   T[  �/��"    A�CNAAA HCA� @   �[  4���`    A�A�C a,D0HA�A�L ��P(E,A0H   @   �[  P���`    A�A�C ^,G0PA�A�D ��P(E,A0H   @   \  l����    A�A�C l,K0VA�A�L ��P(E,A0H      P\  ����       @   d\  �����    A�A�C l,K0VA�A�L ��P(E,A0H      �\  ���       @   �\  �����    A�A�C l,H0bA�A�C ��P(E,A0H       ]  8���       @   ]  D����    A�A�C l,H0bA�A�C ��P(E,A0H      X]  ����       @   l]  �����    A�A�C s,K0VA�A�E ��P(E,A0H      �]  Ȭ��
          �]  Ĭ��       @   �]  Ь���    A�A�C s,H0bA�A�L ��P(E,A0H      ^  ���
          0^  ���           D^  $���Z    A�Cx \A� 0   ^  `����   �#A�BE��h.k
�A�A�C      �^  ���B           �^  X���T    A�A�P�A�x   �^  �����    A�A�A�A�C L
A�A�A�A�IG,G0A4A8A<A@N S,G0A4A8A<A@H CA�A�A�A�4   P_  Ȯ��@    CWBAA HJCBAA H   H   �_  Ю��@    A�A�A�YCEA HBAAA HC�A�A�  D   |_  Į���  �#A�BF���M
�A�A�A�Gd.�
�A�A�A�D   4   `  L���;    A�CMAD HOBAA HA�4   �_  T����   �#A�BF���`.g
�A�A�A�M  T   �`  ����E   A�A�A�A�C@.LIPATCXC\A`L@~
A�A�A�A�L   h   �`  ����   A�A�A�A�C0\
A�A�A�A�Ie
A�A�A�A�Gf<A@ADCHCLAPH0 4   �`  �����   �#A�BF����.L
�A�A�A�A  4   0a  P���  �#A�BF���e.x
�A�A�A�A 4   ha  8���K  �#A�BF����.}
�A�A�A�A  4   �a  P����  $A�BF���e.�
�A�A�A�A L   0b  �����    A�A�A�C p,H0VA�A�A�I ���P(E,A0H       �b  ط��       0   <b  Է���   =$A�BE��h.k
�A�A�C   @   �b  ����@    A�A�CPAD HOBAA HA�A�   4   �b  �����   `$A�BF����.L
�A�A�A�A  4   �b  $���  s$A�BF���^.x
�A�A�A�A 4   $c  ���@  �$A�BF����.}
�A�A�A�A  4   \c  ����  �$A�BF���^.�
�A�A�A�A L   �c  l����    A�A�A�C p,H0VA�A�A�I ���P(E,A0H       <d  ����       0   �c  �����   �$A�BE��h.k
�A�A�C   @   �d  T���@    A�A�CPAD HOBAA HA�A�   4   pd  P���  �$A�BF���.�
�A�A�A�A  4   �d  8���A  %A�BF���e.�
�A�A�A�A 4   �d  P����  %A�BF���.�
�A�A�A�L  4   e  �����  9%A�BF���e.�
�A�A�A�H L   �e  @����    A�A�A�C v,H0zA�A�A�O ���P(E,A0H       �e  ����       0   �e  �����   Y%A�BE��h.k
�A�A�C   @   @f  X���@    A�A�CPAD HOBAA HA�A�      �f  T���{    A�u�    �f  ����           �f  ����1    A�CF eA� D   �f  �����  |%A�BF���E.�
�A�A�A�Cb
�A�A�A�K   4   �f  H���f   �%A�BF���_.P
�A�A�A�AL. 0   Xg  ����]    A�A�C^C HlA�A�  0   �g  ����R    A�CLA VKA HQA�      �g  ����    A�CE LA� (   �g  �����    A�n
�AI
�GJ�   ,   h  8����    A�A�A�|
�A�A�A   @h  ����          Th  ����          hh  ����          |h  ����       H   8h  �����  �%A�BF���f.<
�A�A�A�R`
�A�A�A�MC.   P   �h  �����  �%A�BF���G.E
�A�A�A�HF
�A�A�A�GY
�A�A�A�D $   0i  ����    Cp
MJ
FCE     Xi  ����    CBEE H   xi  ����-    SBEE M   �i  ����       D   Ti  ����c  �%A�BF���z.�
�A�A�A�TD
�A�A�A�AL.  ,   �i  ����6    A�CU
A�FCA LA�L   $j  ����W    A�A�A�C `
A�A�A�GG,A0P KA�A�A�   8   j  �����  &A�BF���|.
�A�A�A�AT.   8   Xj  H����  0&A�BF����.#
�A�A�A�I].  0   �j  ����`    A�A�CG
A�A�ECE  8    k  ����;    A�A�A�`DAA JE�A�A� L   \k  ����v    H�A�A�e
�A�A�OG
�A�A�GCE HGE H   �k  ����          �k  ���          �k  ���          �k   ���          �k  ���          l  ���          $l  ���          8l  ���          Ll  ���          `l  ���          tl  ���           �l  ���$    A�CN LA� X   �l  ����    A�A�A�A�E t
C�A�A�A�MP$A(A,C0H V(A,A0E    0   m  `���?    A�CS
F�CCA ETA� \   <m  l����    A�A�A�A�E {
C�A�A�A�FP$A(A,C0H V,A0E j,A0E  4   Dm  ����q   q&A�BF���t
�A�A�A�PG.   $   �m  $���    A�CLA HC�      �m  ���#    A�R
�MA�   P    n  (���d    A�A�C m
A�A�LC(D,D0A4A8A<A@F<C GA�A�  4   tn  D���X    C e
HC(D,D0D4D8A<A@F<C G   �n  l���"           �n  ����4    A�Q
�NR�   H   �n  �����    A�C^
A�MZ
F�PS
A�LCA EZA E   4   0o  ���c    A�CX
A�Cg
A�HCA E     ho  P���6          |o  |���       $   �o  x���N    A�h
�GK
�EL�$   �o  ����?    CY
DUBA E      �o  ����B    A�Z
�E`�      p  ����          p  ����@          ,p  ���          @p  ���          Tp  ���          hp   ���          |p  ����          �p  ���          �p  ���          �p   ���          �p  ����          �p  ����       <   �p  ���Z    A�CU
A�FZA EL
A�CGA�      4q  $���          Hq   ���          \q  ���E          pq  X���          �q  T���    C$E(D,D0H   �q  T���           �q  P���!    A�CK LA�    �q  \���          �q  h���          r  d���          r  `���2    CZ
CHE    8r  ����          Lr  ����    CS
A     hr  ����          |r  ����          �r  ����          �r  ����          �r  ����          �r  |���          �r  ����          �r  ����          s  ����       $   s  |���!    A�CPA HC�  L   Ds  ����p    A�A�CQ
A�A�H[
A�A�CCA JSBA E L   �s  ����|    A�A�C X
A�A�A[
A�A�CG,A0J W(B,A0E  T   �s  �����    A�A�A�C e
A�A�A�B]
A�A�A�PC$K(A,A0E   @   <t  ���b    A�A�Cb
A�A�GCA J[
A�A�B     �t  8���J    A�CE A� x   �t  d����    A�A�CI HGA HFA HGA HIA HGA HI
A�A�NCH HPK HWA�A�4   �t  �����   }&A�BC���m.F
�A�A�A�C  4   Xu  0���H    A�A�CI FDAA kA�A�0   8u  H���p   �&A�BB��I.L
�A�A�A  �   �u  ����_   A�A�A�A�C@qHBLAPH@PLAPH@JLAPK@sHGLEPFLAHALAPNLAHALAPFLAHBLAPLLAHCLAPH@C
C�A�A�A�IWLAPM@�LAPJ@RHBLAPE@OLAPJ@VHBLAPE@      �v  ���          �v   ���          �v  ���          �v  (���          �v  $���          �v   ���          w  ,���       0   �v  (���J   �&A�BB��P.U
�A�A�E       Tw  D���    A�CE LA� 4    w  @���D   �&A�A�Ea
A�A�ACI       �w  X���.    A�E[ KA�    �w  d���       4   �w  `���*   A�A�C�
A�A�ACB H  4    x  X���*   A�A�C�
A�A�ACB H  0    x  P���B   �&A�BB��V.M
�A�A�E       �x  l���    A�CE LA� 0   Xx  h���B   �&A�BB��V.M
�A�A�E       �x  ����    A�CE LA� <   y  ����^    A�A�CL HZ
C�A�IYC�A�   X   Hy  �����    A�A�A�PA HTC FGA YD
�E�A�LH
�A�A�A       �y  ����.    CQDA FN x   �y  ����N   A�A�A�C0[
C�A�A�JC8D<A@F0A8B<B@BDBHALAPCLC0P<C@F0`
C�A�A�C   p   Dz  ����(   A�A�A�A�C c,C0F B,A0A4C8A<F@H U
A�A�A�A�NO
A�A�A�A�M   �z  `���b   A�A�A�A�C@SLCPF@NLCPF@�DAHALDPH@QDDHCLAPH@R
A�A�A�A�D
A�A�A�A�MCHDLAPF@|DGHALDPATAXD\C`H@`DAHALAPK@]
LEPIQ
LEPJCLAPH@^LAPH@`DAHELCPH@O
LEPEFLCPJ@NDAHGLAPL@P
LEPE�   �{  �����   A�A�A�A�C0�<C@F0R4A8A<A@H0E
C�A�A�A�KS8H<D@F0~4A8A<D@H0E
C�A�A�A�DT4E8A<A@N0Y
C�A�A�A�Ad
<E@E     �|  ����+          �|  ����1    A�o�  @   h|  ���  �&A�BF����
�A�A�A�OD.O
�A�A�A�A   }  ����
       (   }  ����7    A�CT
A�GCC O0   D}  ���`    A�CTA HUA H_A�  <   x}  0���8   A�BF����
�A�A�A�Gr
�A�A�A�A  D   �}  0���[    A�CJ FM
A�NIF C$C(D,A0FIA�   �    ~  H���`   A�A�A�A�F�p�C�F�K�G�A�A�D�A�F�`�D�A�F�^
A�A�A�A�AC�A�E�D�L�g
A�A�A�A�LC�D�A�F�  d   �~  �����    A�A�A�A�C,_0H G
C�A�A�A�EG$A(A,A0J DA�A�A�A� |     ,����   A�A�C d(A,A0M(B,B0A4A8A<A@E<C t$C(A,A0H P
C�A�Cp
C�A�L�$B(E,A0H   �   �  ����   A�A�A�A�CPZ\C`JPE\A`LPuTBXB\A`JP[
A�A�A�A�MF\C`FPgXB\D`AdAhAlApElYPJ
A�A�A�A�D{XE\A`YPIXE\A`LP L   P�  ����    A�A�C,Y0H Q(B,B0D4D8A<A@E<U F
C�A�G   �   ��  X����   A�A�A�C,I0H K,A0H H,A0H J
A�A�A�GX,C0F ],C0F O,C0F M(C,B0B4B8A<A@C<K S
A�A�A�E],A0H C,I0F4A8A<A@K ]$C(A,C0H  $   d�  D���u    A�I
�FV
�J      ��  ����          ��  ����
          ��  ����
          ȁ  ����          ܁  ����
          ��  ����
          �  ����          �  ����
          ,�  |���
           @�  x���K    A�CR sA� D   �  ����  �&A�BF���^.k
�A�A�A�KF
�A�A�A�AY.  $   T�  l���6   'A�CK aA� 4   |�  �����   'A�BF���{.\
�A�A�A�A   4   ��  �����   -'A�BF���e.m
�A�A�A�A  4   �  t����   A'A�BF���p.\
�A�A�A�A   4   $�  �����   U'A�BF���^.m
�A�A�A�A  4   \�  d����   i'A�BF���.N
�A�A�A�A  4   ��  ���  �'A�BF���e.L
�A�A�A�A �   $�  �����    A�A�A�C,L0H M$A(D,A0P K,A0K t
C�A�A�CI(A,B0B4B8A<A@C<C P,A0H RC�A�A�     ��  <���       4   ��  8���\    A�CLFD HX
A�EVA�  4   ��  `���\    A�CLFD HX
A�EVA�  4   0�  ����\    A�CHFD HX
A�IVA�  4   h�  ����\    A�CLGA HX
A�GVA�  4   ��  ����\    A�CLGA HX
A�GVA�  4   ؅   ���\    A�CHDD HX
A�KVA�  @   ��  (���7  �'A�BF���.v
�A�A�A�O^
�A�A�A�A@   ��  $���7  �'A�BF���.x
�A�A�A�M^
�A�A�A�AD   @�   ���V  �'A�BF���e.t
�A�A�A�K^
�A�A�A�A   D   ��  8���V  �'A�BF���e.v
�A�A�A�I^
�A�A�A�A   @   І  P����   (A�BF���p.H
�A�A�A�L^
�A�A�A�A@   �  �����   %(A�BF���p.J
�A�A�A�J^
�A�A�A�A@   X�  �����   <(A�BF���{.H
�A�A�A�A^
�A�A�A�A@   ��  $����   S(A�BF���{.J
�A�A�A�O^
�A�A�A�AD   ��  ����   j(A�BF���^.Y
�A�A�A�M^
�A�A�A�A   D   (�  ����   ~(A�BF���^.[
�A�A�A�K^
�A�A�A�A   D   p�  ����   �(A�BF���e.Y
�A�A�A�F^
�A�A�A�A   D   ��  X���   �(A�BF���e.[
�A�A�A�D^
�A�A�A�A   8   X�  0���=    A�CH HG
A�DEJA HCA�8   ��  4���=    A�CH HG
A�DEJA HCA�8   Љ  8���=    A�CH HG
A�DEJA HCA�$   ��  <���=   �(A�CK hA� ,   ܉  T���[   �(A�A�C` sA�A�,   �  ����[   �(A�A�C` sA�A�$   <�  ����X   �(A�C\ rA�    ��  ����       $   x�  ����X   �(A�C\ rA�    ��   ���       0   ��  ����   �(A�A�Cf WA�A�   $   �  x���a   �(A�C\ {A�    h�  ����       $   $�  ����a   �(A�C\ {A�    ��  ���       $   `�   ���_   �(A�Cc rA�    ��  8���          �  4���       $   ��  0���h   �(A�Cc {A�    0�  x���          D�  t���          X�  ����          l�  |���          ��  x���
          ��  t���          ��  p���       $   ��  |���(    CT
AAADE      �  ����+    C[
ACD    �  ����          �  ����          ,�  ����6          @�  ����6          T�  ���3          h�  0���6          |�  \���6          ��  ����6          ��  ����6          ��  ����	          ̍  ����          ��  ����          �  ����          �  ����          �  ����          0�  ����          D�  ����          X�  ����          l�  ����          ��  ����          ��  ���          ��   ���
          ��  ����
          Ў  ����          �  ����
          ��  ����          �  ����       $    �  ����'    CV
AAAAE      H�  ����          \�  ����       D   p�  ����q    A�CjAAD HC
C�NL
C�AAAEE    ��   ���9    A�e
�J   $   ؏  @���    A�CHA HC�  $    �  8���    A�CHA HC�     (�  0���          <�  ,���          P�  (���       L   d�  $����    A�A�A�A�C0b
A�A�A�A�C]4D8D<A@H0  $   \�  ����   �(CIDAD H 0   ܐ  ����%    A�CE HADAD HA�  H   �  ����T    A�A�A�]
�A�A�NCHAA JJ�A�A�  t   \�  ����}    A�A�A�A�C ]
A�A�A�A�H_$A(A,A0H G
C�A�A�A�ICF�A�A�A�  $   |�  ����   �(CIDAD H 0   ��  ����%    A�CE HADAD HA�      0�  ����A    A�X
�G`�   \   T�  ����j    A�A�F�A�C g$A(E,D0H S
A�A�A�A�DCC�A�A�A�$   \�  ����   �(CIDAD H 0   ܒ  ����%    A�CE HADAD HA�     �  ����       \   $�  ����i    A�A�A�A�C \
F�A�A�A�D\$A(E,A0H GC�A�A�A�$   ,�  ����   �(CIDAD H 0   ��  ����%    A�CE HADAD HA�     ��  ����       \   ��  ����m    A�A�A�A�C0u4A8E<A@H0G
C�A�A�A�HCF�A�A�A�$   ��  ����   �(CIDAD H 0   |�  ����%    A�CE HADAD HA�  (   ��  ����E    A�A�A��A�A�t   ܔ  ����}    A�A�A�A�C ]
A�A�A�A�H\$A(E,A0H G
C�A�A�A�HCF�A�A�A�  $   ��  ���   �(CIDAD H 0   |�  ����%    A�CE HADAD HA�      ��  ����G    A�X
�Gf�   0   ԕ  $���3    A�A�C\AA MA�A�  H   �  0���[    A�A�A�cQAA HF
�A�A�AAAEE   l   T�  D����    A�A�A�A�C0{4P8A<A@SA�A�A�A�A0����A
4A8E<E@EA4A8E<E@   H   Ė  d���=    A�A�A�A�C,N0H$L(A,A0MA�A�A�A�  `   �  X���j    A�A�A�A�C _,D0H$P(D,A0MA�A�A�A�A ����A$A(E,E0D   t�  d���Z    A�A�CcLDA MA�A�A��AAEE    ��  |���          З  x���          �  t���          ��  p���          �  l���           �  h���          4�  d���#          H�  ����       0   \�  |���v    A�CPA RA�A�CE   X   ��  �����    A�A�A�A�H O$D(B,A0H O$D(A,A0H K
C�A�A�A�H   �  ����    CDBB N   �  ����     CDFD N   ,�  ����          @�  ����       4   T�  ����2    A�CP
A�KCAA HCA�      ��  ����#    A�L
�CN�   ,   ��  ����@    A�C T
A�GP(E,A0H  �   ��  ����   A�A�A�A�C@sDEHALAPH@^
A�A�A�A�E�
A�A�A�A�KCDAHALAPL@UDAHALAPL@MDAHALAPH@fHALAPH@  ,   ��  8���5    A�CVBBA JJA�    ��  H���"       0   Ě  d���0    A�A�CTA JEC�A�  0   ��  `���0    A�A�CTA JEC�A�  0   ,�  \���3    A�A�CTA JJA�A�  (   `�  h���(    A�CPA JGA�   (   ��  l���$    A�CPA JCA�   0   ��  p���.    A�A�CVA JCC�A�  @   �  l���@    A�A�C[A JC
C�A�AAAAE    0   0�  h���3    A�A�CTA JJA�A�      d�  t���    CFEBA H D   ��  p���F    A�A�C`AAA HC�A�A��AAEE 8   М  x���4    A�A�A�PBAA JN�A�A� 8   �  |���X    A�C U
A�FN$A(A,D0R NA�   t   H�  �����    A�A�A�A�C h$A(A,A0H P$D(A,A0H C
C�A�A�A�OG
C�A�A�A�AC,E0$   ��  ����"    CJ D$E(B,A0H  ,   �  ����$    A�CJ D$C(B,A0HC� @   �  ����A    A�CYA D$B(A,A0HA�A�AAEE  @   \�  ����=    A�A�A�OH B$B(A,A0JN�A�A�   H   ��  ����_    A�A�A�A�C ~
A�A�A�A�EA$A(E,E0     �  ����&       $    �  ����$    CJ D$B(G,A0H  X   (�    ��O    A�A�A�MDAA HNADA HC
�A�A�AL�A�A�   d   ��  �����    A�A�A�kA A$A(B,A0HA
�A�A�AWAAA JhAAA JSE (   �  L ��    A�CHDA HC�   8   �  @ ��L    A�A�A�q
�A�A�EAAEE  ,   T�  T ��!    A�CE HAAD HA�    ��  T ��       ,   ��  P ��!    A�CE HAAD HA� �   Ƞ  P ��q   A�A�A�A�C s,A0A4B8A<A@H C
A�A�A�A�AN$B(C,A0L T$A(A,A0H E
A�A�A�A�HX
C�A�A�A�BC$A(A,A0H U$A(A,A0H U$A(A,A0H F
$A(E,E0EC,E0   ��  � ��       H   ��  � ��\    A�A�A�A�C {
A�A�A�A�EA$A(E,E0  0   �  ��%    A�CE HAADD HA�      <�  ��    CIADD H 0   `�  ��3    CRBAA HAAAEE      ��  ��       X   ��   ���    A�A�A�GDCG JWAAA JK
�A�A�Mb�A�A�   X   �  T���    A�A�A�A�C@UDKHELAPJ@P
A�A�A�A�EdHALAPH@   4   �  ���B   �(A�BQ
�LF.I
�AM�   X   ��  ����    A�A�A�A�C a(A,A0L M$A(A,A0H L
C�A�A�A�P      ��  ���       d   �  ����    A�A�A�A�C x(A,A0L S$A(A,A0H L
C�A�A�A�Cq$A(E,E0   h   p�  H���    A�A�A�A�C s(A,A0J [
C�A�A�A�IS$A(A,A0H K(C,A0J \,E0    ܤ  ���       ,   �  ���!    A�CE HAAD HA�     �  ���       ,   4�  ���!    A�CE HAAD HA� \   d�  ����    A�A�A�A�C k(A,A0J O$D(A,A0H L
C�A�A�A�Cs,E0 H   ĥ  ���w    A�Ca
A�JDAAA HC
A�MT
A�ECE    �  (��    CBDD HD   0�  (��b    A�A�A�_AA JR
�A�A�NO�A�A� D   x�  P��d    A�A�A�_AA JT
�A�A�LQ�A�A�    ��  x��H       ,   Ԧ  ���X    C a
LC$B(E,A0H I
D L   �  ����    A�A�A�C r
C�A�A�CP(E,A0H E$B(E,A0H    T�  $��       4   �   ��u   )A�BF���c.d
�A�A�A�C   4   H�  h��o   )A�BF���Y.h
�A�A�A�C   0   ��  ���L   $)A�BE��R.N
�A�A�C   p   �  ����    A�A�A�A�C O$F(B,C0H M$A(A,A0H K
C�A�A�A�NS
F�C�A�A�B  x   ��  ����    A�A�A�A�C W
,E0MC$F(B,C0H M$A(A,A0H K
C�A�A�A�AS
F�C�A�A�B D   ��  ���T    A�A�C d$G(A,A0NA�A�A ��A$A(E,E0<   D�  ��?    A�CYAAA HC�C�AAEE    D   ��  ��S    A�A�CfDAA NA�A�A��AAEE x   ̩  ,���    A�A�A�A�C W
,E0MC$F(B,C0H M$A(A,A0H K
C�A�A�A�AS
F�C�A�A�B     H�  P��$    CFDGA N P   �  \���  4)A�BF���W
�A�A�A�M. t
�A�A�A�JU
�A�A�A�H $   ��  ���"    CI A$D(D,D0H  H   �  ���d    A�A�A�A�C C
A�A�A�A�EA$A(E,E0 ,   4�  ���(    A�CE I$D(D,D0HA�    d�  ���       $   x�  ���)    CQ A$G(C,A0H  @   ��  ���3    A�A�A�OA I$G(C,A0HA�A�A�      �  ���%          ��   ��%          �  ��           �  (��%          4�  D��%       4   H�  `��7    A�HKA HDDAA NA�       ��  h��$    CFDGA N    ��  t��          ��  p��           ̬  l��     CBDDD N     �  h��     CBDDD N     �  d��     CBDDD N 0   8�  `��$    A�CP
A�AAAAA H      l�  \��#    CB HKEA      ��  h��#    CB HKEA      ��  t��#    CB HKEA      ح  ���#    CB HKEA  $   ��  ����   H)A�BB��Z.   $   ̭  ����   X)A�BB��Z.   $   ��  \���   h)A�BB��Z.   $   �  ����   x)A�BB��Z.   $   D�  ,	���   �)A�BB��Z.   $   l�  �	���   �)A�BE��I.  $   ��  ,
���   �)A�BB��Z.   $   ��  �
���   �)A�BB��Z.   $   �  �
���   �)A�BB��Z.   $   �  d���   �)A�BB��Z.   $   4�  ���m   �)A�BB��Z.   $   \�  ���   �)A�BF���^. $   ��  ����   *A�BC���c.     �  ��#    CB HKEA  $   Я  ��B   *A�BB��R.      P�  8��           d�  4��!    A�CK LA� 0   0�  @���   (*A�BE��Y.f
�A�A�G   T   d�  ���S  <*A�BF���
�A�A�A�Fz
�A�A�A�Cv.c
�A�A�A�A\.     �  ���          (�  ���           <�  ���!    A�CK LA�    `�  ���           t�  ���!    A�CK LA� \   ��  ����    A�A�A�A�C P,H0D4A8D<A@F X
A�A�A�A�EZ(A,A0J �   ��  `��o   A�A�A�A�C`@hAlApH`!dDhDlApDtAxD|A�U`�hAlApH`O
A�A�A�A�HQ
C�A�A�A�IY
A�A�A�A�A�lMpGtAxD|G�J`blMpGtAxD|G�F`  �   ̲  ���Q   A�A�A�A�C@DDDHDLDPH@]DAHDLAPF@
C�A�A�A�GhHALAPH@]
A�C�A�A�ATA�C�A�A�      d�  ���          x�  ���          ��  ���          ��  ���       <   ��  ���~    A�A�A�r
�A�A�I^
�A�A�P  4   ��  ���|    A�CkD HC
A�A\
A�C     ,�  <��    CP    D�  D��          X�  @��          l�  <��          ��  8��          ��  4��          ��  0��          ��  ,��          д  (��          �  $��          ��   ��          �  ��           �  ��          4�  ��          H�  ��          \�  ��       (   p�  ��I    C\AA HH
OH   ,   ��  ,��X    A�C j$B(D,A0L UA�    ̵  \��          �  h��           ��  d��!    A�CK LA� @   �  p��a    A�A�C`AA HG
C�A�F\C�A� p   \�  ���z    A�A�A�A�C b(A,A0H N
A�A�A�A�KC
F�A�A�A�DTA�A�A�A� P   ж  ����    A�A�CdAA HG
C�A�BSAA Hj
C�A�E     $�  ��          8�   ��           L�  ���!    A�CK LA� 8   �  ��?   �*A�A�CLA HV
A ECA      ��  ��    CF     ķ  ��    C   ط   ��    CF     �  ���          �  ���          �  ���          ,�  ���       0   @�  ���I    C[
BE
ACB HKEA      t�  ��	          ��   ��       0   ��  ���z    A�A�CH HT
D�A�B     и  H��<       (   �  t��m    A�CB HT
C�K      �  ���I       @   $�  ���c    A�HWNA HG
A�ACB HKEA       h�   ��          |�  ��           ��  ��!    A�CK LA�    ��  $��           ȹ   ��!    A�CK LA�    �  ,��    CBEB       �  ,��    CBEB    �   ,�  ,���    A�A�A�A�C@EDAHDLAPATBXA\A`J@u
A�A�A�A�FQ
A�A�A�A�KJLAPDTAXA\A`I@       ��  ���#    CB HKEA      غ  ���#    CB HKEA      ��  ���#    CB HKEA       �  ���#    CB HKEA     D�  ���           X�  ���!    A�CK LA� l   |�  ���:   A�A�A�A�C@MHALAPH@R
A�A�A�A�Lh
C�A�A�A�BkHALAPH@  \   �  ����    A�A�A�A�C0w
A�A�A�A�NV8A<A@H0KF�A�A�A�   \   L�  ���Q    A�A�A�A�C Q$A(A,A0H G
A�A�A�A�B[A�A�A�A�$   T�  ���r  �*A�BE���.     Լ  $��4    CV
G     �  H��          �  D��           �  @��!    A�CK LA� $   <�  L��(    CE HGE HC  8   �  T���  �*A�LB���.I. X.A
�A�A�A   ��  �$��'    CBE \      ��  %��'    CBE \      �  %��       ,   ��  $%��g    A�Cx
A�CV
A�I       $�  d%��<    CLAE MN 4   �  �%��  +A�BF���C.m
�A�A�A�D     ��  h&��       @   ��  d&��P    A�A�C [,A0HA�A�E ��P(E,A0H       ؾ  p&��    A�CE LA� 4   ��  l&��P   ,+A�BF���P.L
�A�A�A�A      4�  �&��          H�  �&���    A���    d�  '���    A���    ��  �'��    CF H  0   ��  �'��A    A�A�CaD KGC�A�     п  �'��    CF H  0   �  �'��A    A�A�CaD KGC�A�      �  �'��     CDD R      @�  �'��          T�  �'��          h�  �'��          |�  �'��           ��  �'��%    A�CO LA�    ��  �'��          ��  �'��          ��  �'��       4   ��  �'���   A+A�BF���@._
�A�A�A�A  4   ��  0(���   Q+A�BF���d.w
�A�A�A�A     `�  �(��<    A�z�  0   $�  �(���   _+A�BB��B._
�A�A�A  4   X�  8)���   o+A�BF���b.x
�A�A�A�A  4   ��  �)���    A�A�C�
A�A�ACB H  0   ��  �*��B   }+A�BB��V.M
�A�A�E       T�  �*��    A�CE LA�    x�  �*��#          ��  �*��           ��  �*��2    A�C\ LA�    ��  �*��          ��  �*��2    A�l�  4   ��  +���   �+A�BF���].L
�A�A�A�A     ,�  \+��          @�  h+��           T�  d+��    A�CL GC�     x�  `+��    A�CL GC�    ��  \+��       P   ��  X+��s    A�A�C\DDA HA�A�L��CA JSBA E      �  �+��2    A�l�  4   ��  �+���   �+A�BF���\.L
�A�A�A�A  �   X�   ,���   A�A�A�A�C0m<A@J0h
A�A�A�A�E�
A�A�A�A�GB<D@H0k<D@H0b<D@H0d<D@H0t<D@H0`<C@F0g<C@F0Y<A@V0 D   ��  8.��k  �+A�BI���[.0n
�A�A�A�H|
�A�A�A�AK.  D   ��  `/��.  �+A�BI���W.0[
�A�A�A�O]
�A�A�A�A.   0   8�  H0��  8,A�BH��m.t
�A�A�B~. 8   l�  $1��0  x,A�BG�A
��A^
��FF.I.  ,   ��  2��  �,A�BG�E
��Av.y. D   ��  3���  �,A�BF���M.�
�A�A�A�Ez
�A�A�A�Am. P   x�  �4��s    A�A�C\DDA HA�A�L��CA JSBA E   8   t�  �4��
  0-A�BI����
�A�A�A�DF.�.   P   �  �6��s    A�A�C^ADA HA�A�M��CA JSBA E   8   �  �6��  d-A�BG�b
��Dd
��LF.G.    8   @�  �7���   �-A�BG�t
��BF.m
��AS.    4   |�  D8���   �-A�BG�b
��DU.n
��A`. 8   ��  �8��:  .A�BG�M.M
��LL
��D_.   4   ��   :��  X.A�BE��b.o
�A�A�Eh.    8   (�  �:��  �.A�BD�X
��AH.q
��A`.    @   d�  �;���   �.A�BG�h.Q
��MI
��Ga
��A`.    <   ��  �<���   /A�BH��x
�A�A�KU. ^
�A�A�C`. 8   ��  H=��  T/A�BF���B
�A�A�A�Bd. M.   8   $�  ,>��  �/A�BF���H
�A�A�A�LT. M.      ��  ?��       D   t�  ?��W  �/A�BC���`.a
�A�A�A�Fi
�A�A�A�D  8   ��  $A��  �/A�BG�[
��Ke
��KF.G.       P�  �A��          d�  �A��          x�  �A��          ��  �A��       P   ��  �A��z    A�A�A�\
�A�A�O\
�A�A�BCA JMBA E    ��  B��          �   B��          �  ,B��G    A�u
�J      <�  \B��          P�  hB��       D   �  tB��  $0A�BI���U.0S
�A�A�A�I]
�A�A�A�A.      ��  LC��       D   h�  HC��  l0A�BI���U.0S
�A�A�A�I]
�A�A�A�A.      �   D��       D   ��  D��  �0A�BI���U.0S
�A�A�A�I]
�A�A�A�A.      d�  �D��       D    �  �D��  �0A�BI���U.0S
�A�A�A�I]
�A�A�A�A.      ��  �E��       D   |�  �E��  D1A�BI���U.0S
�A�A�A�I]
�A�A�A�A.      �  �F��       D   ��  �F��  �1A�BI���U.0S
�A�A�A�I]
�A�A�A�A.      x�  pG��       D   4�  lG��  �1A�BI���U.0S
�A�A�A�I]
�A�A�A�A.      ��  DH��       D   ��  @H��  2A�BI���U.0S
�A�A�A�I]
�A�A�A�A.      0�  I��       D   ��  I��  d2A�BI���U.0S
�A�A�A�I]
�A�A�A�A.      ��  �I��       D   H�  �I��  �2A�BI���U.0S
�A�A�A�I]
�A�A�A�A.      ��  �J��       D   ��  �J��  �2A�BI���U.0S
�A�A�A�I]
�A�A�A�A.      D�  �K��       4   X�  �K��B    A�A�C,a0F,A(A,A0PA�A�L   ��  �K��9    A�A�A�KDA FADA FABA HC�A�A�H   ��  �K��S    A�A�C�A�N0U4A8A<A@H0XA�A�C�A�     ,�  �K��       @   @�  �K��f    A�A�A�}A HM
�A�A�HA�C�A�4   ,�  �K���   <3A�BD�j
��OG.n
��A   4   ��  ,L��Q    A�Cg
C�BCAD HMC�     ��  TL��       $   ��  PL��,   P3A�BH.I
�A   0�  XL��       <   D�  TL��n    A�A�C{A HM
C�A�FIC�A�   ��  �L��       L   ��  �L��Q    A�A�A�A�J b,A0H$A(A,A0H HA�A�A�A�(   ��  �L��$    A�A�CL HE�A�H   �  �L��h    A�A�EKD HP
E�A�LCD HTC�A�   0   �  �L��E   d3A�BB��Z.L
�A�A�A      ��  �L��       P   ��  �L��P    A�A�C\E`F\AXE\A`HPM\A`HPBTBXB\A`JPEC�A� $   ��  �L��    A�CHA HC�     $�  �L��          8�  �L��       @   L�  �L��P    A�A�C [,A0HA�A�E ��P(E,A0H      ��  �L��           ��  �L��!    A�CK LA�    ��  �L��           ��  �L��!    A�CK LA�     �  �L��           �  �L��!    A�CK LA�    8�  �L��           L�  �L��!    A�CK LA�     p�  �L��    A�CE LA� @   ��  �L��P    A�A�C [,A0HA�A�E ��P(E,A0H      ��  �L��           ��  �L��!    A�CK LA�    �  �L��           $�  �L��!    A�CK LA�    H�   M��           \�  �L��!    A�CK LA�     ��  M��    A�CE LA� 0   L�  M��:   u3A�BB��S.L
�A�A�A   $   ��  M��    A�CHA NA�  $    �  M��    A�CHA NA�  $   (�   M��    A�CHA NA�  $   P�  �L��    A�CHA NA�  0    �  �L��:   �3A�BB��S.L
�A�A�A   $   ��  �L��    A�CHA NA�  $   ��  �L��    A�CHA NA�  $   ��  �L��    A�CHA NA�  4   ��  �L��  �3A�BF���Y.�
�A�A�A�C  4   �  �M��$  �3A�BF���Y.�
�A�A�A�C  4   <�  �N��  �3A�BF���h.�
�A�A�A�E  0   ��  �O��4    A�A�MU
A�A�ACE       �  �O��          �  �O��          (�  �O��       4   ��  �O���   �3A�BF���\.Y
�A�A�A�A  ,   t�  P��H   A�C�
A�MCE H     ��  4S��          ��  0S��           ��  ,S��!    A�CK LA�    ��  8S��~    A�GC���(   �  �S��g    A�DB��J
�A�A�M T   <�  �S��   A�A�A�A�C �
A�A�A�A�PS$I(E,A0H Y(A,D0    ��  �T��          ��  �T��           ��  �T��!    A�CK LA�    ��  �T��           ��  �T��!    A�CK LA� 4   ��  �T��o  �3A�BF���L.
�A�A�A�I l   ��  �U��  4A�BF���l.N
�A�A�A�JY
�A�A�A�D^
�A�A�A�OY
�A�A�A�DY
�A�A�A�C   0   ��  �V��T    SE HGE HEEE HH     ��  �V��          �  �V��          �  �V��          0�  �V��*          D�  �V��          X�  �V��          l�  �V��          ��  �V��       ,   ��  �V��)    A�C,H0H$E(A,A0HC� ,   ��  �V��)    A�C,H0H$E(A,A0HC�    ��  �V��           �  �V��!    A�CK LA� H   ,�  �V��Y    A�A�C e
A�A�DG$A(A,A0B,M MA�A�      x�  �V��          ��  �V��          ��  �V��          ��  �V��       8   ��  �V��J    A�C b
A�IC$A(A,A0F,C GA�(   �  ���2    CEEE HEEE H   0�  �V��          D�  �V��          X�  �V��          l�  �V��           ��  �V��!    A�CK LA� <   ��  �V���    F�A�A�C�F
�A�A�A�L`����8   ��  W��F    A�A�A�x
�A�A�CA�C�A� P    �  W��   A�A�C�A�{NR
�C�A�A�JQ
�C�A�A�J 4   t�  �W��[    A�A�Z
�A�COPA
�A�O T   ��  X���   Q�A�A�A�F N
A�A�A�A�D�
A�A�A�A�C  ,   �  �Y��h    C�C�C�_
�A�A�F 0   4�  �Y��o    A�C c
A�HG$M(E,F0Q   8   h�   Z��t    A�A�C�C�E
�A�A�A�P       ��  DZ��S    I�g
�PC�       ��  �Z��?    A�f
�II
�A,   ��  �Z��U    Q�D�y
�A�AC�A�     �  �Z��#       <   0�  �Z���    A�A�A�xBEA HS
�A�A�P  $   p�  �[��}    C�A�O
�A�L     ��  �[��q       4   ��  L\��i    A�A�G|
A�A�IVA�A� `   ��  �\���    A�A�A�^
�A�A�MHADA JL
�A�A�JiAB HXB U  P   H�   ]���    A�A�A�A�G<A@H0I4F8E<A@R0XA�A�A�A�   T   ��  L]���    A�A�A�A�ETAXE\E`PPOTFXE\C`PPbA�A�A�A� <   ��  �]���'   A�BC����
�A�A�A�A�
�A�A�A�A  <  4�  ���.   A�A�A�A�C0H
A�A�A�A�MD4M8E<A@I0t4M8E<A@I0d4M8E<A@I0d4M8E<A@I0s
A�A�A�A�I`4M8E<A@I0�4M8E<A@I0d4M8E<A@I0�4M8E<A@I0c4M8E<A@P0O4M8E<A@P0O4M8E<A@P0O4M8E<A@P0O4M8E<A@P0O4M8E<A@P0O4M8E<A@P0�   t�  ����   A�A�A�A�EP�
A�A�A�A�AC\B`QPI
A�A�A�A�AC\B`QPI
A�A�A�A�AoTMXE\A`PPc
A�A�A�A�ACTMXE\A`PPJTMXE\A`PPPTGXE\E`F\E`HPCTMXE\A`IPQTMXE\A`PP�   l�  �����   A�A�C�A�G0g<F@R0v
A�A�A�A�JQ4F8E<A@P0f<F@R0d4F8L<A@P0Q4F8L<A@P0]4M8E<A@S0z<F@R0H4F8L<A@P0  �   �  ����&   A�A�C�A�G0�4M8E<A@P0Z<T@P0G<S@R0I
A�A�A�A�Fz<a@P0n4M8E<A@S0t4M8E<A@P0O4M8E<A@P0O4M8E<A@P0  �   ��  <���5   A�A�C�G I
A�A�A�H�
A�A�A�PC$F(L,A0P ]$F(L,A0P t$F(L,A0P L$F(L,A0P   @   D�  �����    Q�A�A�C F$M(E,A0I [A�A�A�  p   ��  P���2   A�A�C�A�C0y
A�A�A�A�JG
C�A�A�A�SK4M8J<A@I0g4M8E<A@P0 \   ��  ���`   Q�A�A�A�H �,E0M K
C�A�A�A�Ny
A�A�A�A�C    \�  ����   A�A�A�A�CPh\I`HPM
A�A�A�A�O�
\I`Sd
A�A�A�A�H_\H`OPx
\F`LK
\G`Ft
\H`ZOTHPU
\F`Ig\A`LPE
\H`Xj\C`OPE
\H`mJ
\H`OJ
\F`I�\F`UP�\F`UP�\A`SP�\A`SPR\H`JPB\F`NPC
\F`I|
\F`I�\I`JP�
\I`Ed
\I`E�\I`JP�
\H`iW
\G`I]
\H`EC
\H`E�\H`nPR\I`LPd
\C`E�TAXE\A`HP`\H`_P�
\H`iW
\G`IaTAXE\A`HP`
\H`Zg\A`LPn
\H`VMTAXE\D`HPq\H`nPUTAXE\A`HP`
\H`Z`
\H`\O\H`JPKTAXE\D`HPITAXE\E`HPETAXE\A`HPc\H`JPE\H`]Pz\A`LPg\A`QPu
\H`X�\H`JPx
\A`E~\H`JPH
\F`Ig
\H`OK\I`LPy
\H`Os
\A`E\A`QP_\H`JPQ
\H`LJ
\F`IJ
\H`OJ
\H`O�   l�  ܰ��   A�A�C�A�CP�\A`SP\I`LPp
A�A�A�A�Hd\I`JP�
A�A�A�A�D\H`nPu\H`JP]\F`NPi\I`LP�\H`_Pq\H`JPz\A`QPu
\H`ZJ
\A`Ex
\H`OOTHP  |  D�  $���#   A�A�A�A�E0j
A�A�A�A�I�<H@J0\<H@J0C
A�A�A�A�G�<A@Q0M<H@[0D<H@n0@<A@U0V<H@_0i<H@J0_<I@L0n<A@Q0s<I@J0^
<A@Ep
<A@EL<F@N0�<A@Q0�<A@Q0�<A@S0z
<H@Od<I@J0�<F@R0y<I@N0x<H@J0~<H@J0B<F@N0~<H@J0�4A8E<G@L0t4A8E<A@L0w<F@r0m<I@J0m<I@J0m<I@J0�4A8E<A@L0M4A8E<A@L0E4A8E<E@H0`<H@]0�<H@J0M4A8E<A@H0p4A8E<A@H0o<H@r0P<I@J0W<H@N0l<A@Q04A8E<A@H0I4A8E<A@H0E4A8E<A@H0`<H@a0O
<H@Oa4A8E<A@L0x4A8E<A@L0w<F@t0R<I@L0n<A@U0I4A8E<A@L0M4A8E<A@L0E4A8E<E@H0`<H@_0r4A8E<A@H0p4A8E<A@H0o<H@n0R<I@J0{4A8E<A@H0I4A8E<A@H0E4A8E<A@H0`<H@]0R<I@N0p<H@J0d<H@J0h<F@N0n4A8E<A@L0u<F@r0R<I@J0u
<H@OI4A8E<G@L0M4A8E<A@L0M4A8E<A@L0E4A8E<E@H0`<H@]0A<A@Q0x
<A@Eg<A@Q0Q
<A@EN
<F@Sn
<H@On
<H@Oi<A@S0q
<H@O�<F@N0\<F@N0Q
<H@Oh
<A@EJ
<F@SN
<A@E}
<H@Oa<H@J0@<H@J0
<A@EN<F@N0M<F@T  ��  ����4   A�A�A�A�E@�LAPQ@ELJPN@g
A�A�A�A�GU
A�A�A�A�G@LIPN@p
A�A�A�A�E�LIPN@iLIPN@bLHPJ@eLIPN@YLIPN@YLIPN@GLFPR@gLHPN@�LIPN@ILHPJ@�LAPQ@�LIPJ@�LFPN@bLIPJ@�DAHELAPH@pLHPn@dLHPJ@VDAHELAPH@ADAHELAPH@IDAHELAPH@EDAHELAPH@`LHP]@RLIPJ@jLHPJ@VDAHELAPH@lDAHELAPH@pLHPn@nLAPQ@v
LHPO]LHPJ@[DAHELAPH@IDAHELAPH@EDAHELAPH@`LHP]@RLIPJ@v
LHPOj
LAPEJ
LHPO`LAPQ@_
LAPEkLHPJ@LHPJ@QLHP D   �  �����    A�A�A�A�C0|<I@J0H
A�A�A�A�N4   d�  D���d    A�A�E\H JC
A�A�F   (   ��  |���[    Q�Fo
C�GIA�  p   ��  �����   A�A�A�A�C0
A�A�A�A�Cu<G@O0C
A�A�A�A�NqA�A�A�A�  h   <�  �����   A�A�A�A�E0�
A�A�A�A�CP<H@M0N
C�A�A�A�Gm<H@O0   �   ��  �����   A�A�A�A�E@A
C�A�A�A�PL
C�A�A�A�N
LCPNiLCPO@xLHPS@ILCPJ@/LAPQ@E
C�A�A�A�A�
LAPE    P�  ����$   A�A�A�A�E0�
C�A�A�A�G_
A�A�A�A�M\<H@J0C
A�A�A�A�K�<F@N0O<I@L0S<I@J0f<H@J0W<I@J0w<I@J0e<I@J0O<I@J0O<I@J0~<C@O0e<I@J0s<I@J0O<I@J0U<I@J0U<I@J0O<I@J0O<I@J0O<I@J0j<I@J0  �   t�  ����7   A�A�A�A�C0S
C�A�A�A�Pc<A@Q0�<I@J0�<H@]0g<H@J0R
C�C�A�A�Ec
A�A�A�A�IC
A�A�A�A�I�<H@l0^<H@J0{<A@Q0b<I@J0P
<H@ZJ
<A@E�
<H@Oe<H@J0 <   h�  ���D   A�BC����
�A�A�A�AP
�A�A�A�A �   ��   ���m   A�A�A�A�C0o
A�A�A�A�FU<A@H0K4D8A<A@R0M
C�A�A�A�LT
A�A�A�A�HC<A@L0s<D@H0      @�  ����7    Cd
I  l   \�   ��9   A�A�A�C G
A�A�A�Py
A�A�A�DI
A�A�A�DM
A�A�A�P   h   ��  � ��u   A�A�A�C0}
A�A�A�Jo
A�A�A�Ng
A�A�A�F�
A�A�A�B(   8�   ��A    A�A�C�y�A�A�,   d�  $���	   A�BC����
�A�A�A�A p   ��  ����   A�A�F�A�L`NhAlNpL`Pl\pJ`
A�A�A�A�D�hGlDpS`thGlDpN`   <   �   ���   A�A�C�A�Q��
A�A�A�A�D�   H�  ����   A�A�F�A�S���E�D�L��
A�A�A�A�Nl�G�D�H�M�G�D�H�>
A�A�A�A�A  <   ��  ���D   A�A�F�A�O�'A�A�A�A�  <   �  ���t    A�A�C�S
�D�A�CA
�H�A�F t   T�  4���    A�A�C�A�S�U�C�A�F�B�E�B�E�E
F�A�A�A�LF
F�A�A�A�A  �   ��  |���    A�A�C�H�f�D�A�A�C�B�B�B�I�V�A�A�C�B�B�B�E�q�D�A�A�C�B�B�B�I�P
A�A�A�CF
F�A�A�Bh   |�  ����   A�A�C�A�N@�
A�A�A�A�JY
A�A�A�A�Aj
A�A�A�A�A4   ��    ��X    A�A�Nz
A�A�DEA�A�     �  ( ��       (   4�  $ ��k    A�NB
A�NIA�    `�  h ��          t�  d ��          ��  p ��          ��  l ��          ��  h ��       (   ��  d ��D    A�N(E,H0H K
A�P   ��  � ��          �  � ��       D   �  � ���    A�A�C�K��
C�A�A�AFC�A�A�     `�  !��       D   t�  !��c   A�BD����P��
����PO
����A������� 8   ��  <"���    A�BD����P�O
����A|������ ,   ��  �"���    A�BD����P��������8   (�  @#���    A�BE������
����H}������      d�  �#��    CNAB EC 0   ��  �#���    A�BB��o
�A�A�JI�A�A�   ��  ($��       (   ��  $��A    A�A�C�y�A�A�   ��  <$��       P   �  H$���    A�A�A�C j$C(E,D0I u$O(C,D0I Z
A�A�A�J L   d�  �$���    A�A�A�C m$A(A,D0P a$H(B,A0P HA�A�A�<   ��  %��w    A�Nb
A�NG
F�CS
F�GCC�  0   ��  T%��h    A�NW
A�Ic
C�JFA�P   (  �%��/   A�A�C�A�N@\
C�A�A�A�J�C�A�A�A� D   |  l&��{    A�A�A�C [(I,H0H,A(M,K0dA�A�A� X   �  �&��   A�A�D�P,A0H Y
A�A�A�En(A,F0P Q
A�A�A�G  T     X'��f   A�A�A�E@�HDLAPY@K
A�A�A�Es
F�A�A�A   <   x p(��'   A�A�C�C@�HJLAP]@AA�A�A�\   � `)��I   A�A�A�G0�8J<A@L<A8J<A@S0|
C�A�A�ICC�A�A�   D    P*���    A�A�A�C g(E,A0f,A(E,A0fA�A�A� �   ` �*��n   A�A�C�A�N`�
A�A�A�A�P�lCpH`�hDlApNlAhDlApP`WlHpL`MlHpL`qlFpL`�dBhClApI`SlIpH`C
A�A�A�A�AwhJlHpNlAhDlApR`�lCp]`ndDhDlDpI`~lDpH`klGpT`ylHpH`    \ 1��V    A�T�    x P1��W       0   � �1��c    A�A�NMB d]A�A�     � �1��K          � 2��K           � P2��V    A�NB CA�P    �2���    A�A�N t
A�A�Jc
C�A�IF,E0L G
A�A�A     ` (3��       (   t $3��2    A�NMA PCA�   H   � 83��    A�A�A�A�N0v8E<D@T0F
C�A�A�A�A    � 4��            �3��%    A�Ba�       4��    A�BU�     @ �3��    A�BV�     ` �3��%    A�Ba�     � �3��    A�B[�     � �3��    A�BW�     � �3��+    A�Bg�     � �3��"    A�B^�        4��    A�B[�       �3��     A�B\�     @ �3��     A�B\�     ` �3��!    A�B]�     �  4��=    A�By�     � 4��;    A�Bw�     � 84��    A�B      � '4��    A�BV�     � !4��     A�B\�      !4��!    A�B]�     < "4��!    A�B]�     \ #4��=    A�By�     | @4��    A�BT�     � 84��+    A�Bg�     � C4��1    A�Bm�      � T4��    A�BA�K�A�      A4��&    A�Bb�       G4��y    A�Bu�    @ �4��4    A�Bp�     ` �4��;    A�Bw�     � �4��     A�B\�     � �4��     A�B\�     � �4��     A�B\�     � �4��     A�B\�      	 �4��;    A�Bw�      	 �4��8    A�Bt�     @	 5��     A�B\�     `	 5��8    A�Bt�     �	 5��    A�BX�     �	 5��    A�BX�     �	 5��    A�BA�     �	 �4��
    A�BF�      
 �4���    A�B      
 H5��.    A�Bj�     <
 V5��    A�BI�     \
 C5��U    A�BQ�    |
 x5��Q    A�BM�    �
 �5��S    A�BO�    �
 �5��   A�B��    �
 �6���    A�B�� (   �
 /7���   A�BE��s�A�A�       ( �9��e   A�BD�]��   L �;���   A�B��   l G=��R   A�BN�    � y>��   A�BD���A�   � Z?��J    A�BF� $   � �?��A   A�BG�5�A�       � �G��c   A�BG�X��     �L���	   A�BD��	��   @ �V��i    A�Be�    ` �V��C   A�B?�$   � Y���   A�BG���A�   $   � �e���   A�BG���A�   $   � 4n���   A�BD���A�   (   � �r��   A�BE���A�A�       $ �x���   A�BG����   H U����    A�B��     h �����   A�BG����   � O����   A�B��   � ����   A�B��   � �����   A�B��   � p����   A�B��    )���J   A�BF�   , S���8    A�Bt�     L k����    A�B��    l 3���4    A�Bp�     � G���D    A�B@�    � k���*    A�Bf�     � u���#    A�B_�     � x���    A�BZ�      v����    A�B��    , ���
    A�BF�     L Л��
    A�BF�     l ����     A�B\�     � ����V    A�BR�    � ���!    A�B[�     � ���    A�BT�     � ���    A�BU�      ���\    A�BX�    , ���    A�BN�     L ���,    A�Bh�     l ���9    A�Bu�     � 5���5    A�Bq�     � J����    A�B��    � ����b    A�B^�    � �����    A�B��     ����q    A�Bm�    , ܝ��    A�B{�     L ;���j   A�BD�b��   p ����
    A�BF�     � k���o    A�Bk�    � ����|    A�Bx�    � ���)    A�Be�     � ���8    A�Bt�       7���K   A�BD�C��   4 ^���A    A�B}�     T ���;    A�Bw�     t ����I   A�BE�   � ã��    A�BX�     � ����G    A�BC�    � ���W    A�BS�    � ���    A�BR�      ���6    A�Br�     4 )���F    A�BB�    T O���;    A�Bw�     t j���J   A�BF�   � ����5    A�Bq�     � ����1    A�Bm�     � ����Y    A�BU�    � ���    A�BT�      ���    A�BH�     4 צ���    A�B��    T y���8    A�Bt�     t ����U    A�BQ�    � Ƨ��;    A�Bw�     � ����    A�B��    � ����)    A�Be�     � ����%    A�Ba�      è���    A�B��    4 ����e    A�Ba�    T ũ��    A�BU�     t ����     A�B\�     � ����     A�B\�     � ����    A�BR�     � ����    A�B[�     � �����    A�B��     ���+    A�Bg�     4 $���    A�BV�     T ���    A�B[�     t ���8    A�Bt�     � 5���;    A�Bw�     � P���     A�B\�     � P���X    A�BT�    � �����    A�B��     ����`    A�B\�    4 5���    A�BW�     T 0���    A�B      p )���    A�B      � +����    A�B��    � ����v   A�Br�   � ���3    A�Bo�     � ���3    A�Bo�      ���=    A�By�     , 6���p    A�Bl�    L ����B    A�B~�     l �����    A�B��    � ���2    A�Bn�     � -���c    A�B_�    � p���%    A�Ba�     � u���1    A�Bm�      ����
    A�BF�     , p���'    A�Bc�     L w���*    A�Bf�     l ����#    A�B_�     � ����:    A�Bv�     � ����    A�BZ�     � ����Y    A�BU�    � հ���    A�B��     ^����    A�B��    , ̱��@    A�B|�     L ���    A�BR�     l ����    A�B��    � P����    A�B��    � �����    A�B��    � W���    A�BA�     � <���    A�B        0���u   A�BD�m��    , �����   A�BD����    P ����{   A�BD�s��   t S���     A�B\�     � S���c    A�B_�    � ����[    A�BW�     � ѷ���    A�BD���� ,   � v���%   A�BI����A�A�A�      ( k���]    A�BY�    H ����I    A�BE�    h ����    A�BU�     � ����    A�BV�     � ����    A�BU�     � ����    A�BV�     � ����"    A�B^�      ����%    A�Ba�     ( ����     A�B      D ����    A�B      ` ����"    A�B^�     � ����"    A�B^�     � ����    A�BU�     � ����    A�BV�     � ����    A�BW�       ����?    A�B{�       ����-    A�Bi�     @ ����T    A�BP�    ` ���3    A�Bo�     � #���0    A�Bl�     � 3���-    A�Bi�     � @���T    A�BP�    � t���    A�BT�       l���6    A�Br�       ����-    A�Bi�     @ ����T    A�BP�    ` ����    A�BV�      ��&4  f,� �� �  �� �� ��  ��'�  �� �� �  �� �� �4  ��&� 5� eK  ��Y  n�� �  ��L  �� �&     � ��  ��	��          � (-S"u �  �/u         � 	    �	 ��	\l �   � 9(QB  q� �  �� �� �  �   }       @	� 5%Ux�� �  �� �� �  �   }      @	� 9*T�w  �� �  �� �� �  �   }     @	� 9)Dqg  �� �  �� �� �  �   }      @	��	[k �     � A0  ;�X� �B  �  �� �� �� ��  }       @	� =.�  ���� �� �  �� �� ��  }     @	� 9*  5!�9  �� �� �� �  ��  }     @	� E4�  ����  �o��� �� �� �  ��  }       @	� E7  d��� �x  �H��� �  �� �� ��  }    @	� E7  d��� �x  �H��� �  �� �� ��  }    @	� E7  y��� �s  �H��� �  �� �� ��  }    @	� E7  p��� �|  �H��� �  �� �� ��  }    @	� E7  p��� �|  �H��� �  �� �� ��  }    @	� E7  j��� �r  �H��� �  �� �� ��  }    @	� E7  j��� �r  �H��� �  �� �� ��  }    @	� E7  d��� �x  �H��� �  �� �� ��  }    @	� M?�  ������������ �  �� �� �   }    @	� M<'  ���  ���  ���� �  �� �� �   }       @	� I6  T��)  �
8��
�
�� �  �� �� �   } }       @	� M=1  j�������
��� �  �� �  �� �   } }    @	� M=+  _���������� �  �� �  �� �   }      @	��+ &  9  ��+ &  9  ��7Z U  h  ��  1� �  ��+ &  9  ��3   A  ��3   A    � )  � ;� x��=��  ��       ��*9 G  ��)8 F  ��,; I  ��*9 G  ��)8 F  ��,; I  ��+� |� �  �  ��+� |� �  �  ��(7 E  ��'6 D  ��)8 F  ��)� |� �  �  ��0? M  ��/> L  � K�r� �  ��      ��+ 9  ��+ 9  ��  Wu �  ��  Wu �  ��+ 9  ��� g� �  �    � �u  >,�
��
��
�(�
���������������������
��
���	�
�
� �    }     � ��  �(�������������������������������������	��	��	��	��
��
"  �� �    }      � ��  �(�������������������������������������	��	��	��	��
��
"  �� �    }      � ME/  ��� ��� �
;� �����  � � �� �  �� �       � ME/  ��� ��� �
;� �����  � � �� �  �� �       ��(P� ��� �     � -"��  �����  �� �          � )!E�  �����  �� �       � -"��  �����  �� �          � -"��  �����  �� �          � -"��  �����  �� �          � %E����  �� �         � %E����  �� �         � %E����  �� �         ��  ]� u�� �  ��  ]� u�� �  ��
9s� �  ��  H�� �  ��(  ��� ��  �� ��  �i� �  ���� �  ���� �  ���� �  ���  ��� ��  ���  ��	� ��  ���  ��� ��  ���  ��� ��  ���  ��	� ��  ���  ��
� ��  ��D ?  R  ��,�� �� �� �� �  �  �  �    � +MZ        ���}� �  �  ��< @ h  ��  ]� �  ��  &<� �  ��0� ?� j� y� �� �  ����� �  ��i� �� �  ��/  �� �  ��n� �� �  ��/  �� �� �� �  ��n� �� �� �� �  ��0� ?� j� y� �� �  ��$  �� �  ��g� �� �  ��$  �� �� �� �  ��g� �� �� �� �  ��0� ?� j� y� �� �  ��,  H� �� �#  ��n� �� �  �� ,  H� �� �� �� �  ��n� �� �� �� �  ��0� ?� j� y� �� �  � N��  �� �   �	� (<HOX            ��o�� �  � P�\��&    }    � )C��������               � E���� �       � =2f  ������������ �  �          ��W^ l  ��3 [� �  ��N] k  ��1 ,  E  ��+ ?  ��/ *  =  ��/ *  =  ���� �    � )'�z  �� �� �   }     @	�� ��/  Dd Tf �  ��n� �� �  ��$  9Y I[   ��g� �� �  ��,  H� z� �� �(  ��n� �� �� �  ��,  H� z� �]� �(  ��,  H� z� �]� �(  ��n� �� �Y� �  ��n� �� �Y� �  ��$  9� I^� �  ��$  9� I^� �  ��/  D� TS� �  ��/  D� Tc� �  ��g� �_� �  ��g� �_� �  ��n� �X� �  ��n� �X� �  �� �� �� �� �� �� �� �� �� �� �� �� �� �� �� ��   � &0      ��,V p  ��"P j  ��  - G  ��TP  �� ��  ��Z (m K"  ��Z (m K"  ��Z (m K"  ��Z (m K"  ��Z (m K"  ��2  Q� Z� }"  ��Z (m K"  ��Z (m K"  ��Z (m K"  ��Z (m K"  ��Z K"  ��'o 1� `"  ��)s 2� d"  ��/ *  ��  !o �     � A2)�  ���  �$��� �  �� �� �   }     @	� 	1     }         � )FL  ���&  �"� �?   }     �	� IA�9����S���������������  �    }   ��?  L� �   � )B    }    ��.  Il ~  ��
m� �  ��+  Gi {  ��
k� �  ��/ *  =  ��	fv �  ��	eu �   � E5  g��  ���� �  �� �� �  �   }      @	� E5  c��  ���� �  �� �� �  �   }      @	� =.  8�^  �� �  �� �� �  �   }     @	� 1!�  ���� �� �  �   }      @	� 9+.  ���� �  �� �� �  �   }    @	� E5"  V��  ���� �  �� �� �  �   }      @	� 1"�  ����� �� �  �   }     @	� =/  f��  �� �  �� �� �  �   }    @	� 1#  F�d0  �� �� �  �   }    @	� =-  Ete  �� �  �� �� �  �   }      @	� =/  W2��  �� �  �� �� �  �   }    @	� =/$  j��  �� �  �� �� �  �   }    @	� =/   h��  �� �  �� �� �  �   }    @	� =.  2�p  �� �  �� �� �  �   }     @	� 9*"  e��� �  �� �� �  �   }     @	� =/  t��  �� �  �� �� �  �   }    @	� =/!  t��  �� �  �� �� �  �   }    @	��&� ��   � =/  f��  �� �  �� �� �  �   }    @	� E5  a��  ���� �  �� �� �  �   }      @	� E5  a��  ���� �  �� �� �  �   }      @	� E5  a��  ���� �  �� �� �  �   }      @	� E5  a��  ���� �  �� �� �  �   }      @	� E5  a��  ���� �  �� �� �  �   }      @	� E5  a��  ���� �  �� �� �  �   }      @	� E5  a��  ���� �  �� �� �  �   }      @	� E5  a��  ���� �  �� �� �  �   }      @	� E5  a��  ���� �  �� �� �  �   }      @	� E5  a��  ���� �  �� �� �  �   }      @	� E5  a��  ���� �  �� �� �  �   }      @	� Gv        �         � .7     ��' 5  ��' 5     � 
".��          � 
"��          � 
1��          � 
%4��       ��U#� �E� �  ��5�� �  ����{�9���6�����    ����                                                ����   �		�		�		         
	
	
	
	
	
	
	
	!
	%
	)
	-
	
	1
	�P�� 	"	�!	�]@b�fGCC: (GNU) 4.9.1              ��           \    {
       �@   0�K   ��  ���    �s   ��p   �   ��   ��               �+       �*           ,    �,        �P   p�c   ��V               �4       @�E           �   B       ��   ��   ��   М+    �   �%   @��   Н   �    �    �   @�V   ���   p��   `��   `��   P�%   ���   �e   ��a   �T  P�i  ��B  �    �s   ��   ��   Шz   P�   p�   ��G   �    �    �    �   @�   `�   ��R   �R   @�R   ��  ��   ��@    �   �   �   0�   @�   P�  p�   ��  ��   ��  к   �  �    �    �  0�   @�  P�           �    ��       ��   `�   ��$   ��   ��    ��?   0�   @�j   ��   ��M    �I   p��    �    �s   ��Z    �           <    �%      �   ��   ��   �X  ��          �   ΃      ��   ��   ��   ��   ��   ��   ��   �    �   0�   @�   `�   ��   ��   ��   ��   ��   ��   ��   ��    �!   0�   @�   P�   `�   p�   ��   ��   ��   ��   ��&   ��&    �&   P�&   ��&   ��&   ��&   �&   @�&   p�&   ��&   ��m   @�m   ��Z   �   0�   P�!   ��!   ��!   ��!   �   0�!   `�!   ��!   ��   ��!   �!   @�!   p�!   ��"   ��>   �   0�   @�!   p�>   ��m    �   @�   P�!   ��2   ��'  ��@   0�>   p�F   ��F   ��  ���   ���    �(  P�L   ��K   ��N   @�"   p�"   ��S    �S   `�S   ��S    �"   P�H   ��H   ��L   @�K   ��N   ��"   �"   @�S   ��S    �S   `�S   ��"   ��H   @�H   ���    ��   ���   ���   P�   p�>   ��>   ��   �@   P�8   ��J   ��I   0�K   ��"   ��"   ��S   @�S   ��S    �S   `��   0�   P�8   ��8   ��8   �8   P�8   ��   ��4   ��6   0�:   p�2   ��R   �Q   p��   P�   p�   ��   ��   ��   ��G   0 G   � �   �   ��  P   p>   �   �   �    8   @8   �8   �8    8   @   `>   �>   �   �    ,   0   @   P   `�   ��   �>   �.   �    $   0   @�   �L   @	�      X  �L   �L    L   pM  �L   L   `L   ��  @ L   � �   (L   p(L   �(L   )�  �*L    +L   P+L   �+I   �+I   @,I   �,I   �,I   0-I   �-I   �-I    .I   p.I   �.I   /I   `/I   �/�  `1�    25   @2  `:  �B�  `Dw   �D4   G/   PG�    H  K�   N1   @Nr   �N�  `Q1   �Qp   Rr   �R  �S(  �V5    Wo   �W�  PZ5   �Zo    [(  0\(  `]�   `^�  @a7   �a�  `d;   �dc   e�    f  i�  m  0o�   r=  @  `�  ���  0��  ���   Н�  ���
  ��k  �k  `�k  Ю�  ��7   �|   `�d  м�  ��7   ��|   p��  0�7   p�|   ���  ��7   ��l   `�|   ���	  ��7    �|   ���	  P�7   ��|   ���           D    /�      �    �   0�   @�   P�   `�           T    �      ��   ��   p�W   ��   ��"   ��"    �    ��           4    �0      ���  ��%   ��_   P�F          T    T      ��m   �   0�l   ��   ���   p��    �
   0�
               Y�      @�          �   ��      `�6   ��F   ��W   ��"   P�`   ��`   ��   ��   ���   0�   P��   ��   ���   p�   ���    
        @ �   � 
   �     Z   `�   PB   �T    �   �@   �@   0�   ;   @�    E  p	  �
�   p  �K  ��  p�   �    �   �@   0�       @  `�  ��   p   ��   p@   �  �A   �  ��  ��   0   @�   0@           T    ]P      p{   �    1   P �   "f   p"]   �"R   0#           $    ��      P#�   �#�           �    ~�      p$   �$   �$   �$   �$�  @'�  �(�   �)   �)-   �)   �)c  P+6   �+W   �+�  �-�   0`   �0;   �0v   @1           �   �      `1   p1   �1   �1   �1   �1   �1   �1    2   2   02$   `2�    3?   @3�   4q   �4   �4#   �4d   P5X   �5"   �54    6�   �6c   P76   �7   �7N   �7?   08B   �8   �8@   �8   �8   �8    9   9   09   @9   P9   `9   p9   �9Z   �9    :   :E   `:   p:              k      ��   ��   �:   �:!   �:   �:    ;   ;2   P;   p;   �;   �;   �;   �;   �;   �;    <   <    <   0<!   `<p   �<|   P=�   �=b   P>J   �>�   p?�    @H   p@p   �@_          l    ʷ      @C   `C   pC   �C   �C   �C   �C   �CJ   0D   PDD   �D.           L    )�      �D   �D*  F*  @GB   �G   �GB    H           �   $       H^   �H�    I.   0IN  �J(  �Kb   P�   S+   0S1   pS  �T
   �T7   �T`   @U8  �V[   �V`  @X�   �X�  �Z  �\�   �]�  @_u   �_   �_
   �_
   �_    `
   `
    `   0`
   @`
   P`K   �`  �a6   �a�   �b�   Pc�   �c�   �d�   �e  �f�   �g   �g\   �g\   Ph\   �h\   i\   pi\   �i7  k7  PlV  �mV  o�   �o�   �p�   �q�   �r   �s   �t    v    w=   `w=   �w=   �w=    x[   �x[   �xX   @y   PyX   �y   �y�   Pza   �z   �za   @{   P{_   �{   �{   �{h   @|   P|           �   #�      p|   �|   �|
   �|   �|   �|(    }+   0}   P}   p}6   �}6   �}3   0~6   p~6   �~6   �~6   0	   @   P   `   �   �   �   �   �   �   �   0�   @�
   P�
   `�   p�
   ��   ��   ��'   Ѐ   ��   ��q   p�9   ��   Ё   ��    �   �    ��   ��   �%   @�T   ��}    �   @�%   p�A   ��j   0�   P�%   ��   ��i    �    �%   P�   `�m   І   ��%    �E   p�}   ��   �%   @�G   ��3   Ј[   0��   ��=    �j   p�Z   Њ   ��   ��    �   �    �   0�#   `�   p�v   ���   p�   ��    ��   ��   Ќ2   �#   @�@   ���  P�5   ��"   ��0   ��0    �3   `�(   ��$   ��.   �@   0�3   p�   ��F   ��4    �X   ���   �"   @�$   p�A   ��=    �_   `�&   ��$   ��O   ��   Е   �L   @�!   p�   ��!   ��q  0�   P�\   ��%   ��    �3   @�   `��   ��   ��B   К�   p�   ���   P��    �   0�!   `�   p�!   ���   P�w   О   �b   `�d   ПH    �X   ���   �    �u   ��o   �L   `��   ��   ��T   �?   0�S   ���   0�$   `��   �"   0�d   ��(   Ч   �)    �3   `�%   ��%   ��   �%   �%   @�7   ��$   ��   ��   Щ    �    �            �    <�      0�$   `�#   ��#   ��#   �#    ��   ���   @��   Ь�   `��   ��   ���   @��   Я�   `��   �m   `��    ��   ��#   вB           ,    �	       �   0�!   `��               �C	      �S          ,    9b	      p�   ��   ��!           <    �c	      ��   ж!    ��   �o  `�Q              v	      ��           $    �v	      ��   ��           4    S�	      ��    �~   ��|    �           d    ��	       �   0�   @�   P�   `�   p�   ��   ��   ��   ��           D    ��	      ��   ��   ��   ��    �   �I           L    a�	      `�X   ��   ��   ��!    �a   ��z   ��           ,    x�	      ��   ��   ��!           T    T�	      �?   P�   `�   p�   ��   ��   ��   ��           ,    /�	      ��I   �	    �           4    Ƚ	      0�z   ��<   ��m   `�I               ��	      ��c           ,    ��	       �   0�   @�!           $    ��	      p�   ��!           $    �	      ��   ��               <�	      ���           4    ��	      ��#   �#   @�#   p�#           <    =�	      ��   ��!   ��:   ��   ��Q               ]
                  N
      �r              
      ��4               [
              ,    L 
      ��   ��   ��!           T    $
       �(   P��  0�'   `�'   ��   ��g    �<   `�          4    #~
      ��   ��P   ��    �P           L    P�
      P�   `��    ��   ��   ��A   �   0�A           $    R�
      ��    ��               $�
              t    G�
      ��   ��   ��    �%   0�   @�   P�   `��   ���   ��<    ��   ���           ,           P��   P�B   ��           D   6D      ��   ��#   ��    �2   @�   P�2   ���    �   @�   P�   p�   ��   ��s    �2   `��   ���  ��k  @�.  p�  ��0  ��  ���  ��s   �
   �s   ��  ���   ���   ��:  ��   �   ��    ��    �  @�  `�   p�W  �   �   �           z   �   �   �G   0   P   p  �   �  �   �  �          0  P	   `	  �
   �
  �   �  �   �        @   P  p           $    �      �B   �9           �    *B      S   p   �f   ��   �Q   �   �,       0n   �   �Q   $   @h   �E       P               �a      `           �    �      �   �   �P   �    !   0   @!   p   �!   �   �!   �   P   `   p!   �   �!   �   �!       @:   �   �   �   �    :   @   `   �           L    ��      �  �$  �  4   P   `   p           $          ��    H          ,    L<      p!   �!   �!!           ,    K      �!~   @"g   �"          T    �]      �#   �#   �#!   $    $!   P$o  �%  �&T           �    |�      @'   P'   `'   �'*   �'   �'   �'   �'   �')    ()   P(   `(!   �(Y   �(    )   )    )   0)J   ��2           $    ��      �)   �)           ,    ��      �)   �)   �)!               ��      �)�              |�      �9              ��      P�u              ��      ���(              R      �          w
       -
  �  k              �  (  _� �>   �  �  P   �  �  o  �	  �  qW  !~   int   "�   �  #  s  NE   �  VE   .  <s   `  D~   �  Ws   �  _�   �  e~   t   m~   a  u~     ~~   �  �~   3  �~   �  �~   H  �~   y  �~     �~   s  �~   T   �~   �  �~   F  �~   �  �~   �  �~     �~   V  �~   %   �  \	  2~   o  7~   �  <~   �  C~   �  ~   *    �  ~    	rem ~    +   �  #@  A  �  $,    	rem %,    A  &  
std 
 �  	v  	wA  	{�  	�   	�'  	�<  	�Q  	��  	��  	��  	��  	�  	�.  	�N  	�o  	�z  	��  	��  	��  	��   � �~   �  �   �  �  >       �� "  %   �  H~   <     �  I,   Q     �  �   z  z  z  3   3   �   �  �  ~   �  z  z   div   �  ~   ~        ��  �     �   A  �  ,   ,    �  .~       3    �  \3   !  !    3    '    3  >~   N  !    3    �  o  �   3   3   �   k� q~   �  |�  l      W  �    �   �    f,   �    �  ~    �  g>   �    �  ~    ?  �~   �     �  ,1  ��   �8  ptr ,�   � �m
  � �   D  OD   �   �  PD  1  QD  �  Wm   �   ^  Xm  U  =�   �   �   >�  B  ?�  �  E�   �   B   F�  C  G�  e  H�  8  I�  �  J�  

  X    �   �  Y   �
  Z   �   `)  �   �  f:   �   �  g:  �  h:  �  nc   �   �	  oc  �  pc  H  v�   �   `  w�  w  x�     y�  ~  �        ��  �  ��    ��  �   ��  �  ��  �	  ��  �  �       �    �  �  �  �  �O     �  �O  �  �O  �  �O  m  ��   $  	  ��  2	  ��  �  ��  9  ��  [  ��   /  J  ��  �  ��  7  ��  �  ��   :  I	  ��  $	  ��  �   �#   E  N  �#  p  �@   P  �  �@  :  �@  �  �@  d   �@  �  Ɂ   [    ʁ  �  ˁ  �	  Ѫ   f  �  Ҫ    ��   q  �  ��  �  ��  �  ��  +  ��   |  �  ��  �   ��    �%	   �  �
  �%	  �  �%	    �N	   �     �N	  F  �N	  �  �w	   �  �  �w	  �  �w	  �  3�	   �  �  4�	  �   8�	   �  �  9�	  l	  =�	  �  N  >�	  ^  ?�	  L  @�	  a  D
  �  B  E
  �	  F
    G
    H
  y  I
  �   \
   �  �  !\
    ;�     x!   �  �  �  k  (      �  �  (  _� �>   �  �  P   �  �  o  �	  �  qW  !~   int   "�   �  #  s  NE   �  VE   .  <s   `  D~   �  Ws   �  _�   �  e~   t   m~   a  u~     ~~   �  �~   3  �~   �  �~   H  �~   y  �~     �~   s  �~   T   �~   �  �~   F  �~   �  �~   �  �~     �~   V  �~   %   �  \	  	2~   o  	7~   �  	<~   �  	C~   �  
~   *    �  ~    	rem ~    +   �  #@  A  �  $,    	rem %,    A  &  
std  R  v  wA  {R  �n  ��  ��  ��  �	  �$  �9  �T  �o  ��  ��  ��  ��  ��  �  �8  �W  � �� Zg  �� Wg  �  ��   �� ?  k    �z ;  �z L4  <    �  r  �  f.   � �~   g  g   m  �  >�  �  �   �� �  %   �  H~   �  �   �  I,   �  �   �  �   �  �  �  3   3   �   �  �  ~   	  �  �   div   $  ~   ~        ��  9  �   �   A  T  ,   ,    �  .~   o  �  3    �  \3   �  �  �  3    �    3  >~   �  �  �  3    �  �  �   3   3   �   k� q~   �  |�  l      W�    �     �    f,   8  �    ~    �  g>   W  �    ~    ?  �~   l  �      3  A  P>  �  A]	   t  Bn	  +  F�  �  G�  �  Jt	  p  N~   p  Y~     Zz	  �  [z	   �  \\  $w  ]�   (4  a�  0 =  Pp�    s�    �  xn	  +  |�  �  }�  �  �t	  p  �~   p  �~     �z	  �  �z	   �  �\  $w  ��   (4  ��  0 �  ��  �  �t	   �  �l    W  `3  �  r   �  �
    �   �  }�     �   �  �t	  ,  �   �  W3  B  r   �  �t	  W  �    �  ��   m  t	   8  ^�  �  ~   /	  r  �  :	     ��  �     P  @X    ++CCUNG }  LX   ++CCUNG�  ��  �   !�  [  "�  �:    �   #�  r�  o�   !  �    $�  ��  �    �  %abi �l  + 0l     1~   (  5l   h  7l   �  =�   &B�  �  '�   '�  'M  '3  '�  ']  'K  '	  '�   �  L}  �  W�  �  (�  �  �   �  ^   Z/	  �  \r   �  ]�  V  bF  `  cF   �  n~   @	  )�  *�  ,   *2  >   �  (n	  �    c	  w  �	  P   + l  �  %�	  =  '\   ;  (\  l  )\  -  *z	  w  +z	  �  ,P     -P    C  ��  ,�  
  -c `r     ,�  )
  .exc ��   ,  ?
  -eo }�   ,  U
  .exc ��   /�  �
  0�  �  0�� :	  0�  �   0n  ~   0Q  z	  0�  \  0�  z	  12xh t	    3j  �z	    .p �z	  .val �  14�� �l   4  �P   4�T  �Q	    Q	  5  :3  T  0�� :T  0  :Q  12e <z	  2tmp =Q	    �	  �  6  ~     7    �  8h  �   k  ,,  �  -c Wr   /=  *�  0�  *�  0n  +�  0Q  ,�  0�  -  12xh /t	    �  6~   �  6z	  	  6\  ,B  %  .ptr ͞    ,W  <  0m  �t	     7(  P  Z  8h  Z   <  9�  �z	  �@   ��  :p �z	      :val ��     ;��7   <�� �l   J   <  �P   �   <�T  �Q	  �     E	  =@  �3  0�K   �1  >�  �1  �   >�  �1    >�  �7  0  ;<�8   ?�  ۞   �l  �  �   9�  �z	  ��  ��  >�� �P   \  >WC  �\  �  :p �z	  V  @val ��  � A   n  Bu å  /  �  n  <�T  �g  �  C �   �  Dtmp �E	  �\E�_  FPv FR�\  C0�    M  Gtmp �Q	  H�
  0�    �I�
  J�
  �  ;0�    K�
    K�
  0  K�
  O     A0   d  Ba �g  b   Le�w    M  �Nptr ��   Nu2 �^   Nu4 �l   Nu8 ��   Ns2 �e   Ns4 �~   Ns8 ��     \  3V  Hl   �  O�� HP    9�  [1  ���   �Z  >�� [T  �  :i [Q	  �  PH   Dptr ]\  �lQ�  ��`   _O  J�  >  L��w    LВ=    9�  �3   �s   �^  >�� �T  g  >�  �^  �  >�  �   �  R  �E	  � Px   Be �z	  (  P�   <�  �1  ;  Btmp �Q	  N  S�
  @�'   �1  T�
  �O   J�
  l  ;@�'   K�
  �  K�
  �  K�
      Ur��  E  FPw  E}��  FRu FQ�\    �	  9l  e\  ��p   ��  >�� eP   ,  >�� e:	  M  Lœ~   L�w   L���   L	��    5q  z	     0�� :	  0�� P   -p z	  -val �   9Z  1z	  �  �h  >�� 1:	  �  :p 1z	  �  >�� 2T  ^  P�   Btmp 4Q	  }  <�  5P   �  Q�  G��   <�  J�  �  J�  		  J�  	  J�  F	  US�d  �  FPu FRw  Ee�=  FPu FQv   S�
  ��   I  I�
  J�
  Y	  ;��   K�
  l	  K�
  �	  K�
  �	    Q�
  ���   R]  J�
  �	  J�
  �	  P�   K�
  �	  K�
  
  K�
  &
    L.��     Vm   ��  ��  W�� ^~   � W�  _/	  �W�  `r  �W�  a�  �W�� b:	  �X  vY  Q�Y4  ���A  �  Z�  k�  9
  [�� m�	  �HZQ  nz	  �
  Z�  oz	  �
  \p pz	  �  Z�  q\  �  \ip q\  e  Zn  r~   �  [�  s�   ��Z$� t3  �  [�  u~   ��2xh �t	  ]�  `�8  ��  J�      ^�  ��   �  J�  8  J�  `  J�  �  J�  �  ;��   _�    AP  �  [�  �\  ��[  �\  �@[�  �\  �DZ  �Q	  �  ]�  ��x  ��  J�    J�  S  J�  f  J�  �  U��d  �  FPu FR0 E��=  FPu FQs   ]�  ���  �#  J�  �  J�  5  J�  S  J�  r  UҖd    FPs FR0 E�=  FPs FQu   ]�  ��  ��  J�  �  J�  "  J�  K  J�  j  U��d  t  FPs FR0 E�=  FPs   `�
  ��  �I�
  J�
  �  P�  K�
  �  K�
  "  K�
  n     A�  R  [w  E	  �@[�  E	  �DZ�  1  �  Z�  ^  �  Z�  3  �  Ze  3    ^)
  �   3K  J3
  2   ^  �-   \�  J#  F  J/  [  ;�-   K<  z  KF  �  a�
  ��"   ?J�
  �  J�
  �  ;��"   K�
  �  K�
    K�
  (      U��_  �  FPw FR�@ UƘ_  
  FPv FR�D UD��    FP�H U]��  9  FRu FQ�� E�Z  FP�HFR��  ^U
  v�*   ��  Jn
  G  I�
  I�
  J�
  [  I�
  Jz
  p  Jb
  �  ;v�*   _�
    Lڕ�   L��   L���   L9��   U\�   �  FP�FR��FQ�H Uo�d    FR� L��!  L���  Lҗ;  L%�F  U��   L  FP�FR��FQ�H U��d  a  FR� U��d  v  FR� L�#!  L�F   b�  e'   '}  '�  '�    V�   ��   �  W0  ��   � C,��     Zo  ��  �  c�  �V  d�      Z  `  �   e�  �&  5  8h  /  Z   f�  �B  8h  /  8#  f    gD  ��  [�� ��	  �H2xh �t	  Z�  �z	  �  [�  �Q  V[#  ��  WA  �  Z�  �  �  Z'  �t	    g�  ��   gQ    ^%  ]�   �!  J/    a)
  ]�   �J3
      ^B  њ   	?  JP  *   L[��  Ux�   h  FP0FRuDFQuP U��Z  �  FPuPFQs  L��6!  U��Z  �  FPuPFQ0 LΚ;!  L�N!  L��   ^5  ��   �  IB  L��   L2�  LM�!  LV�#!  L��g!   L��l!   �    6�  hD  O/   �   h�  P/  h1  Q/  h�  WX   �   h^  XX  hU  =u   �   h�   >u  hB  ?u  h�  E�   �   hB   F�  hC  G�  he  H�  h8  I�  h�  J�  h

  X�   �   h�  Y�  h�
  Z�  i�   `  �   h�  f%   �   h�  g%  h�  h%  h�  nN   �   h�	  oN  h�  pN  hH  vw   �   h`  ww  hw  xw  h   yw  h~  �     h   ��  h�  ��  h  ��  h�   ��  h�  ��  h�	  ��  h�  �     h  �  h  �  h�  �  h�  �:     h�  �:  h�  �:  h�  �:  hm  �o   $  h	  �o  h2	  �o  h�  �o  h9  �o  h[  ��   /  hJ  ��  h�  ��  h7  ��  h�  ��   :  hI	  ��  h$	  ��  h�   �   E  hN  �  hp  �+   P  h�  �+  h:  �+  h�  �+  hd   �+  h�  �l   [  h  �l  h�  �l  h�	  ѕ   f  h�  ҕ  h  ز   q  h�  ٲ  h�  ڲ  h�  ۲  h+  ��   |  h�  ��  h�   ��  h  �   �  h�
  �  h�  �  h  �9   �  h   �9  hF  �9  h�  �b   �  h�  �b  h�  �b  h�  	3�   �  h�  	4�  h�   	8�   �  h�  	9�  hl	  	=�  �  hN  	>�  h^  	?�  hL  	@�  ha  	D�  �  hB  	E�  h�	  	F�  h  	G�  h  	H�  hy  	I�  h�  
 G    �  h�  
!G   r  j�   ++CCUNGj�  ++CCUNGkf� ��  �\  �   :	   #  �\  �   :	   )  �\  �   :	   $  ��   :	  ~   F   �  ��   :	  \   �  ��   !  :	     �\  !  :	  !   ~   l�  �   6!  �    m�  l�  �   N!  >    n�  g!  �   �   n	   m�  o>  Y  �     �    _  .  �  k  x      y  std  <   _� ��    �  �  �   �*   ��   sz 0   � ���   ��   ��    �  	�  ��  �   �   
0    >  Y  �   
�      
�            >  k  �      U  std 
 E  v  6�  x  K�  �  ME   x  Ob   m   G  E   	�  Qw  �   �   G   	�  R  �   �   G   
  T8  E  �   �   M   x  Z�   �   G   x  \�   �   G  S   x  _�     G  �   x  c  #  G  ^   �  p�  d  ;  F  G  S   �  t�  d  ^  i  G  ^   �  {y  �  G  j   n	 ~%  �  �  G  d   �  ��  q  �  �  M   �  �h  x  �  M    ;    :;   �  �Y  � �  3�  �� Z�  �� W�  /  m      a�    �  f.   ;   �  �  �  ;   ;   int �  �  (  �  �  �  �  ��   �  ��   #  �� 
  ��  + 0�  �  (  5�  �  =�  �   B�  @  !�   !�  !M  !3  !�  !]  !K  !	  !�   �  L�  �  WV  \  "l  @  l   r  #^   Z�  �  \�   �  ]K  V  b�  `  c�   �  	 j    
 |  #A  P>b  �  A�   t  B�  +  F  �  G  �  J�  p  Nj  p  Yj    Z�  �  [�   �  \�  $w  ]E  (4  ar  0 #[  `d�    g�   $exc i�   #�  ��  �  ��   �  ��   %�  ��  �  l   %�  ��  �  E   &�  Wq  �  �   '�  <  E  �  �   (�  [)P  @�   ++CCUNG)}  L�  ++CCUNG*�  �:  K     +  c]  E   ,�  X<  -�  oE  E    .abi ��  �  "�  E   �  �  /�  �  �  �  0�  b  1�  �  2exc �l   3�     4,�  @  2exc  l  56e  #�    1�  '  2ptr �E   1�  <  7c W�   8�   �P   ��  9�  � 9�  �:�  w  ;  <p�6   =�  >�  =  >�  Q  =�  ;  ?V�K     @�  p�c   �<  Aobj <E  � BU  <�  �B�  =�  �Cx�[   D�  A<  p  6e  E�  <}�]  <��  <��*  <ƛ�  <Λi  <ӛ9    �  @  ��V   ��  C�R   D�  ]<  �  De  ^�  �  E'  �   f�  >1  �   <�]  <��  <$�i  <,�9    �  F   ++CCUNGF"  ++CCUNGG�  �@  �  l   H�  �@  l    L   �  0  �  k  �      �
  �  (  _� �>   �  �  P   �  �  o  �	  �  qW  !~   int   "�   �  #  s  NE   �  VE   .  <s   `  D~   �  Ws   �  _�   �  e~   t   m~   a  u~     ~~   �  �~   3  �~   �  �~   H  �~   y  �~     �~   s  �~   T   �~   �  �~   F  �~   �  �~   �  �~     �~   V  �~   %   �  \	  2~   o  7~   �  <~   �  C~   �  ~   	*    �  	~    	rem 	~    +  	 �  	#@  A  �  	$,    	rem 	%,    A  	&  
std  
  
v  
wA  
{
  
�&  
�M  
�b  
�w  
��  
��  
��  
�  
�'  
�T  
�t  
��  
��  
��  
��  
��  
�  � �� Z  �� W  �  f.   � 	�~        %  �  	>;  ;  B   �� H  %   �  	H~   b  B   �  	I,   w  B   �  	�   �  �  �  3   3   �   �  �  ~   �  �  �   div 	  �  ~   ~        	��  �  B   �  	 A    ,   ,    �  	.~   '  B  3    �  	\3   G  G  B  3    M    3  	>~   t  G  B  3    �  	�  �   3   3   �   k� 	q~   �  	|�  l      	W;  �  B  �   �    	f,   �  B  �  ~    �  	g>     B  �  ~    ?  	�~   $  B   + 0l   (  5l   �  =�   B�  �  �   �  M  3  �  ]  K  	  �   �  LE  �  W�  �  �  �  �   �  ^   Z�  �  \:   �  ]�  V  b$  `  c$        A  P>�  �  A-   t  B>  +  F�  �  G�  �  JD  p  N~   p  Y~     ZJ  �  [J   �  \/  $w  ]�   (4  a�  0 �  W  �  :   �  �D  �  �    P  @0   ++CCUNG }  L0  ++CCUNG!�  �:    �   "�  o�   �     �  #abi ��  �  >  �    3    P  P   $�  %�  q  &c W:   %�  �  'exc Դ   (�  '@�E   ��  )�  '�  � *\  U�   1�  +f  �   ,r�   �  -xh 3D  .}��   .U�  .���   /D  O   �   /�  P  /1  Q  /�  W0   �   /^  X0  /U  =M   �   /�   >M  /B  ?M  /�  Ev   �   /B   Fv  /C  Gv  /e  Hv  /8  Iv  /�  Jv  /

  X�   �   /�  Y�  /�
  Z�  0�   `�  �   /�  f�   �   /�  g�  /�  h�  /�  n&	   �   /�	  o&	  /�  p&	  /H  vO	   �   /`  wO	  /w  xO	  /   yO	  /~  �	     /   ��	  /�  ��	  /  ��	  /�   ��	  /�  ��	  /�	  ��	  /�  ��	     /  ��	  /  ��	  /�  ��	  /�  �
     /�  �
  /�  �
  /�  �
  /m  �G
   $  /	  �G
  /2	  �G
  /�  �G
  /9  �G
  /[  ��
   /  /J  ��
  /�  ��
  /7  ��
  /�  ��
   :  /I	  ��
  /$	  ��
  /�   ��
   E  /N  ��
  /p  �   P  /�  �  /:  �  /�  �  /d   �  /�  �D   [  /  �D  /�  �D  /�	  �m   f  /�  �m  /  ؊   q  /�  ي  /�  ڊ  /�  ۊ  /+  �   |  /�  �  /�   �  /  ��   �  /�
  ��  /�  ��  /  �   �  /   �  /F  �  /�  �:   �  /�  �:  /�  �:  /�  3c   �  /�  4c  /�   8�   �  /�  9�  /l	  =�  �  /N  >�  /^  ?�  /L  @�  /a  D�  �  /B  E�  /�	  F�  /  G�  /  H�  /y  I�  /�      �  /�  !  :  1�   ++CCUNG1�  ++CCUNG ��   �  �C  �L  �V  �      	  �  �� �� (  �  �  �  Z   �  �  o  �	  �  qW  !�   int   "%   #  .  <}   `  D�   �  W}   �  _�   �  e�   t   m�   a  u�     ~�   �  ��   3  ��   �  ��   H  ��   y  ��     ��   s  ��   T   Ȉ   �  Ј   F  ׈   �  ��   �  �     �   V  �   H   �  s  NO   �  VO   \	  2�   o  7�   �  <�   �  C�   �  �   �  �  H   	pO qO !  
std % �:  @	  %+  \%  0a1  vr  �J  N  T  
G   �#  &  _Tp �.  �?  �    �=  	�P  �b  	�H   Fe  	�   �#  	�P  �&  	��  �3  	�=  �  �<  �<   ~  eq 	�<-  �<  �  �<  �<   lt 	��1  �<    �<  �<   ��  	eF  �   '  �<  �<  �   �K  	�9  �  A  �<   �(  	
!  �<  e  �<  �  �<   1  	�A  �<  �  �<  �<  �   �5  	�'  �<  �  �<  �<  �   �3  	�A  �<  �  �<  �  ~   +  	:  ~  �  �<   �  �C  	 �P  �  
  �<   �B  	$6  �<  )  �<  �<   eof 	(�:  �  ?  	,N0  �  �<    E  �[  9Q  p�  G0  s�   �T  t	  %  {�  �  �?   %  ��  �  �?  �   �:  �b;  �  �  �  �?   �T  �4>  �  �  �?  	   �T  �QM  	      �?   �F  ��?  �?  #  .  �?  �    I  �O  �?  F  Q  �?  �   (*  �	H  [  i  t  �?  �   �O  �eT  [  �  �  �?  �   �O  ́?  �  �  �  �?  �?   �$  	   �:  Z�   _� �A   5�<  6�=  7>  �?  �:   K  \z  �:    �e  _�   �4  c*>   �J  d0>  ��  qA  G  H>   ��  sW  b  H>  N>   !W  yn  H>  �     �  �J  p  "�B  �  #�   $%  �   %�B  �  �  e>  �  N>   &�B  �  e>  �      �e  y  '[V  �  �  $�G  !�    <  x�   �4  {   �J  |%   �J  M<   `S  �R<   ~J  �   �J  �  �%  ��  �K  ��   I  ��  :!  �>   %H  �D	  #_   (�3  2�  (�G  7�  (t3  B�>  )�'  ��O  }>  *V  ��N  �<  �  �  �>   *3  �o+  �<      �>   +�P  ��O    %  w>   +�M  ��P  8  >  w>   +�,  �-  Q  \  w>  �   *�+  ��R  �  s  y  w>   *3  �   �  �  �  w>  N>  N>   �/  !�B  w>  �  �  �  N>   +�O  �|6  �  �  w>  N>   ,(  ��6  �  	  w>  N>   -�   �-  �  	  	  w>   .�1  o�*  �  3	  w>  N>  �    -�A  $n%  �  \	  b	  k>   -�A  (�I  �  z	  �	  q>  �   -"A  ,�%  w>  �	  �	  k>   -�1  2E)  /  �	  �	  k>   -�/  6;&  /  �	  �	  k>   ,�>  :�>  �	  �	  q>   -S  A:2  �  
  !
  k>  �  �   ,�#  K�(  5
  J
  k>  �  �  �   -9  S>$  �  b
  r
  k>  �  �   --U  [�7  �<  �
  �
  k>  �   /�5  d�-  �
  �  �  �   /	1  m�P  �
  �  �  �   /�3  v\-  �
  �  �  H    /nU  ��-    �  /  /   /nU  �nG  5  �  ;  ;   /nU  ��   U  �  �  �   /nU  �IP  u  �  �  �   �J  �rR  �   �  �  �   ,�=  ��H  �  �  q>  �  �  �   ,V  �)  �  �  q>   0�'  �D*  }>  1�0  ��  �  q>   2�0  �    q>  N>   �0  �)  4  q>  �>   �0  �D  Y  q>  �>  �  �   �0  �i  �  q>  �>  �  �  N>   �0  ��  �  q>  �  �  N>   �0  ��  �  q>  �  N>   �0  ��  �  q>  �  H   N>   1�0  "�  	  q>  �    3�  *,Q  �>  "  -  q>  �>   3�  2�G  �>  F  Q  q>  �   3�  =�%  �>  j  u  q>  H    3S� f�&  /  �  �  q>   3S� q�>  ;  �  �  k>   4end y<  /  �  �  q>   4end �6;  ;  �  �  k>   3I ��$  S  
    q>   3I ��7  G  )  /  k>   3��  �lC  S  H  N  q>   3��  �CM  G  g  m  k>   3r ��R  �  �  �  k>   3�K  �r5  �  �  �  k>   3�3  �j=  �  �  �  k>   5�� �  �  �  q>  �  H    5�� ��F      q>  �   3I  v  �  (  .  k>   5�E  �|U  C  N  q>  �   5�1  -�  c  i  q>   3�� 5�?  �<  �  �  k>   3�:  D�6  #  �  �  k>  �   3�:  UW    �  �  q>  �   4at k
/  #  �  �  k>  �   4at ��7        q>  �   3�F  ��/  �>  /  :  q>  �>   3�F  �k:  �>  S  ^  q>  �   3�F  ��H  �>  w  �  q>  H    3@  DA:  �>  �  �  q>  �>   3@  U�1  �>  �  �  q>  �>  �  �   3@  )�D  �>  �  �  q>  �  �   3@  ��*  �>    !  q>  �   3@  �6  �>  :  J  q>  �  H    5�G  -aN  _  j  q>  H    �3  �b*  �>  �  �  q>  �>   3�3  ^ 2  �>  �  �  q>  �>  �  �   3�3  �=  �>  �  �  q>  �  �   3�3  z�T  �>  �    q>  �   3�3  � @  �>  !  1  q>  �  H    5� ��E  F  [  q>  /  �  H    3� �\+  �>  t  �  q>  �  �>   3� �u>  �>  �  �  q>  �  �>  �  �   3� g|=  �>  �  �  q>  �  �  �   3� "�@  �>  �    q>  �  �   3� 9k<  �>  '  <  q>  �  �  H    3� K�'  /  U  e  q>  /  H    3bL  d�R  �>  ~  �  q>  �  �   3bL  t�2  /  �  �  q>  /   3bL  �L&  /  �  �  q>  /  /   3�%  �9F  �>  �  	  q>  �  �  �>   3�%  �|<  �>  "  A  q>  �  �  �>  �  �   3�%  ��T  �>  Z  t  q>  �  �  �  �   3�%  ��A  �>  �  �  q>  �  �  �   3�%  b>  �>  �  �  q>  �  �  �  H    3�%  3%  �>  �    q>  /  /  �>   3�%  'V7  �>    6  q>  /  /  �  �   3�%  <�+  �>  O  d  q>  /  /  �   3�%  Q'S  �>  }  �  q>  /  /  �  H    3�%  vj.  �>  �  �  q>  /  /  �  �   3�%  ��9  �>  �  �  q>  /  /  �  �   3�%  �C  �>    0  q>  /  /  /  /   3�%  �>/  �>  I  c  q>  /  /  ;  ;   -�?  ��&  �>  {  �  q>  �  �  �  H    -�1  �O  �>  �  �  q>  �  �  �  �   ,)  �z-  �  �  �  H   N>   6+E  �3J  �    �  H   N>   3�5  ��)  �  '  <  k>  �  �  �   5n	 @D  Q  \  q>  �>   3W�  �6  �  u  {  k>   3�A  %�A  �  �  �  k>   3��  ,Z5    �  �  k>   3�(  �;  �  �  �  k>  �  �  �   3�(  I�%  �       k>  �>  �   3�(  X�5  �  )  9  k>  �  �   3�(  �^   �  R  b  k>  H   �   3�(  v�S  �  {  �  k>  �>  �   3�(  	K  �  �  �  k>  �  �  �   3�(  �o?  �  �  �  k>  �  �   3�(  J5  �  �    k>  H   �   3NW  ��Q  �  $  4  k>  �>  �   3NW  /�I  �  M  b  k>  �  �  �   3NW  ��,  �  {  �  k>  �  �   3NW  ��;  �  �  �  k>  H   �   3�S  ��I  �  �  �  k>  �>  �   3�S  >T?  �  �    k>  �  �  �   3�S  05  �  $  4  k>  �  �   3�S  $S:  �  M  ]  k>  H   �   3�>  2hL  �  v  �  k>  �>  �   3�>  SUB  �  �  �  k>  �  �  �   3�>  Q�2  �  �  �  k>  �  �   3�>  _�K  �  �    k>  H   �   3�4  qT  �    /  k>  �>  �   3�4  j�K  �  H  ]  k>  �  �  �   3�4  ��5  �  v  �  k>  �  �   3�4  N.  �  �  �  k>  H   �   3U+  �)    �  �  k>  �  �   3��  �!1  �   �  �  k>  �>   3��  ��T  �     *  k>  �  �  �>   3��  ��O  �   C  b  k>  �  �  �>  �  �   3��  �;.  �   {  �  k>  �   3��  ��B  �   �  �  k>  �  �  �   3��  ��,  �   �  �  k>  �  �  �  �   �  !T  H   7�E  r  7�F  �   8�&  8�7    �o  >�"   �| C�   9Q  b<   #  9�F c<  9�R  d<  93  e<  9�  f<  9�K  g<  9�@  h<   :all i<  ?;�� ��  $:!  �>   $NF  ��>  $�E  ��  $p0  ��>  $�%  ��>  <S  ��>  <�R  ��>  <3  ��>  <�$  ��>  <�K  ��>  <�@  ��>  <�@  ��>  ,�4  �Z  S  Y  �>   ,�=  y)  m  s  �>   %�� �  �  �>  ?  �   %�� �  �  �>  �  �   %�� �  �  �>  �   %N  �  �  �>  �    %�� �    �>  ?   ,�  �U    #  �>  ?   -�&  �.  �<  ;  A  �>   ,�F  &�;  U  e  �>  ?  #   ,�9  )�Q  y  �  �>  ?  ?   ,WR  ,`2  �  �  �>  ?  �>   ,�S  /=  �  �  �>  �>  �>   =e  7,  �  �>  �>  �    $�$  �>   <OD  �>  <gP  �>  <�F  $�>  >< E   ?< r9   �K  �    @id ��   $�U  ��   <�I  �>  ,�  �<?     �   �>  �>   Aid ��   �   �>  �>   Bid ��   �   �>   C4H  ��(  �  �   �>    �o  u�   �   �>   �o  ~�   !  �>  �>   2�o  �!  "!  �>  �   �o  �2!  G!  �>  �>  �  #   �o  �W!  l!  �>  �>  �>  #   5  �|!  �!  �>  �    �  ��*  �>  �!  �!  �>  �>   H�  ��N  �"  �!  �!  �>   U  �9  �<  �!  �!  �>  �>   2  �t*  �<  "  "  �>  �>   DjP  �D    )"  �>   ERD  �Q  �>  F�o  7J"  U"  �>  �>   G�K  :�N  G�A  =�5  �K  @I  #  �"  #   ,�,  CH<  �"  �"  �>  �>  �>  #   E   #   �     � >  HW  3_#  I�4  I�$  Iq-  Ic=  Io'  I�5   I�%  � I�8  �IX)  �I�%  �I�  �IaO  �IY=  � IP  �� I�C  ��IwS  �I�O  � I�?  �I�5  �� H
$ g�#  I)W  I�   I�U  I�A  I�8  I�P   IEH  �� H�4  ��#  IO   I�7  I(  I�Q  IG  �� H��  ��#  I�R   I�-  I�1  IlO  �� >b4 �&   �P  ��"  J�N  ��#  J�  J�#  3n4 '�T  �#  4$  :$  %C   3�/ v2  3  S$  ^$  �C  3   3l6 ��K  3  w$  }$  %C   3l6 �6N  3  �$  �$  �C  3   3s0 B?  �#  �$  �$  �C  �#   3s0 S�(  �#  �$  �$  �C  �#  �#   J�9  i_#  3*H  ��7  �>  %  %  %C   �#  K�4  %  Ldec %  Kt-  %  Lhex %  Kr'  %  K< %   Loct %  @K� %  �M[)  %   M�%  "%   M�  &%   MdO  )%   M\=  ,%   M�P  /%    M�C  3%   @KzS  6%  �K�O  9%  JM�?  <%  K�7  N1&  $  K(  Q1&  K�Q  V1&  KO  Y1&   Lin wm&  �$  Lout zm&  Lcur ��&  $   �#  N�8  �:�&  �,  ;�_ �$'  $�M  ��<   $N  �?  2�_ .�&  �&  *?  $?   1�.  ��&  '  *?  �    C�  ��3  �<  '  0?    �&  O]-  <"P�  A?    �b  >H    Fe  ?�   �#  @�   �&  A�   {'  ER/   �!  F]-   �E  G�&   '<  I�0  2�  T�'  �'  Q?  �   W?  ]?   Q�@  ]�&  �'  �'  Q?  �   W?   RT  luB  c?  (  (  Q?  i?   RT  u�H  c?  '(  2(  Q?  ~?   RT  �-  c?  J(  U(  Q?  �?   RT  �/  c?  m(  x(  Q?  :    RT  � /  c?  �(  �(  Q?  A    RT  ��.  c?  �(  �(  Q?  �<   RT  [*/  $?  �(  �(  Q?  o    RT  �4/  c?  �(  )  Q?  h    RT  i�Q  $?  )  ')  Q?  �    RT  ��Q  c?  ?)  J)  Q?  v    RT  Ʉ/  c?  b)  m)  Q?  �    RT  ͎/  c?  �)  �)  Q?  %    RT  ��.  c?  �)  �)  Q?  3    RT  ��.  c?  �)  �)  Q?  �<   RT  ��.  c?  �)  �)  Q?  ,    RT  �d9  c?  *  *  Q?  �   RT  w�  $?  4*  ?*  Q?  ]?   Rput ��V  $?  W*  b*  Q?  B'   5�9  7MN  w*  �*  Q?  �?  3   B'  �9  �A  $?  �*  �*  Q?  �  3   � �qP  $?  �*  �*  Q?   �A  �yC  Z'  �*  �*  Q?   3A  E  $?  	+  +  Q?  Z'   3A  !0W  $?  -+  =+  Q?  f'  $   1�  �N+  ^+  Q?  �   W?   Z'  N'  �5  ?�"  $?  �+  �+  ]T  :   Q?  :    �'  sN  ?�$  $?  �+  �+  ]T  A   Q?  A    70  ?�6  $?  �+  �+  ]T  �<  Q?  �<   ;  ?�*  $?  ,  ,  ]T  �   Q?  �    0@  ?�,  $?  >,  I,  ]T  %   Q?  %    6<  ?C;  $?  j,  u,  ]T  3   Q?  3    �S  ?�<  $?  �,  �,  ]T  ,   Q?  ,    =  ?�#  $?  �,  �,  ]T  �  Q?  �   !T  H   7�E  r   �� 
8�,  oS  
8�#    �� 
V-  oS  
V�#    i� 
t+-  TC  
t�     x� 
�D-  V  
��     2� 
�]-  V  
׈     >�E  R/  33F  ;�S  @  -  �-  $@   4tie !�G  Q?  �-  �-  $@   9U  ؍0  $  �-  �-  $@   �M  ��B  $  �-  �-  $@   S`V  ]-  �-  .  .A  �    1aV  �.  .  .A   eU  ��4  ,.  7.  .A  $   bU  �IQ  K.  V.  .A  $   �=  �93  �<  n.  t.  $@   Z  �4O  �<  �.  �.  $@   3[F l�L  �.  �.  �.  $@    �b  KH   3��  ��$  �.  �.  �.  $@  H    3[F ��@  �.  �.  /  .A  �.   !T  H   7�E  r  i3 ~P4  +/  6/  .A  @   T�1  )�%  F/  .A  $    >�M  �0  3�-  �  �@  t/  z/  �@    �b  �H   3�-  P  �@  �/  �/  �@   5� !4  �/  �/  @  �    3�S  �YH  �/  �/  �/  @  z/    Fe  ��  3�W  �B  3  0  0  @  �D  3   z/  3X'  F6  �   <0  B0  @   -9  ��<  o0  Z0  o0  @  {0  $  �$    �#  ��   �&  ��  3:H  ?,  o0  �0  �0  @  o0  �$   !T  H   7�E  r   >"(  �2  4put 	&"  �0  �0  �0  -I  �0  ?  1  :    J�B  �@3  J�b  �H   4put #	z"  �0  21  L1  -I  �0  ?  1  A    4put �F!  �0  e1  1  -I  �0  ?  1  �<   4put )	�"  �0  �1  �1  -I  �0  ?  1  �    4put -	;#  �0  �1  �1  -I  �0  ?  1  %    4put ^	�!  �0  �1  2  -I  �0  ?  1  3    4put b	/K  �0  12  K2  -I  �0  ?  1  ,    4put w	=I  �0  d2  ~2  -I  �0  ?  1  �   !T  H   7QJ  @3   >�+  3  3��  a�)  �2  �2  �2  =D  H    J�b  �H   UKC  3�T  �2  �2  �2  �2  =D  H    =+3  ��3  3  =D    �>  b�  [  `'  
�@3  �>  
�H    !T  H    ;G  ؙ4  5    }'  �R/  (T  ��?   �U  �<   �E  �&  "  ��3  �3  �?  �?   "  ��3  �3  �?  �?   �  �'V  �?  �3  �3  �?  H    3*  )A  �?  �3  �3  �?   3�F  	j8  �?  4  4  �?  �    3�F  �8  �?  84  >4  �?   3V  �0  �<  W4  ]4  �?   3�E  L  �?  v4  �4  �?  �  3   !T  H   �E  r   @3  V0T  �4  %��  :�4  �4  �M  �   !T  H    ]-  R/  W*  K�"  �4  �"  �"   W�*  O�"  
5  �"  �"   W�*  ��#  $5  �#  �#   W*  ��#  >5  �#  �#   W	W  ��B  X5  �B  �#   �#  W	W  [HC  w5  NC  �"   �"  W+  W�"  �5  �"   WwA  _HC  �5  NC  �"   �2  3  W�;  �3  �5  !T  H   �E  r  @  @   XJ  ,6  !T  H   �E  r  $?  �  3   W�   خ<  16  �$  	  �?  �?   WN  .�G  O6  �R  �2  =D   Yp9  J$?  w6  !T  H   �E  r  $?   XG  9�6  !T  H   �E  r  $?  3   Y5  �$?  �6  �E  r  $?  H    Y5  $?  �6  �E  r  $?  �   W�2  .'I  7  �R  �0  -I   �0  >�N  �7  3\�  �DU  �"  ,7  27  "M   3��  �  Q7  K7  Q7  "M   J7# p  3�p  �kV  Q7  w7  }7  "M   3�{  �w:  �7  �7  �7  "M   J�b  oH   3]�  ��H  �7  �7  �7  "M   Zid >E   !T  H    
7  Wf3  p@3  8  !T  H   @3  �  �    ZJ  4�>  $?  78  !T  H   �E  r  $?   �'  @�=  $?  c8  !T  H   �E  r  $?   6�+  
��)  $?  �8  !T  H   �E  r  $?  3   6�+  
m�/  $?  �8  !T  H   �E  r  $?  �,   6�+  
OqM  $?  �8  !T  H   �E  r  $?  �,   6�+  
��:  $?  #9  !T  H   �E  r  $?  -   6�+  
�R@  $?  S9  !T  H   �E  r  $?  +-   6�+  
�R  $?  �9  !T  H   �E  r  $?  D-   6�V  L�L  $?  �9  !T  H   �E  r  $?  �  3   5  �Q$  $?  �9  �E  r  $?  Z    5  ��#  $?  :  �E  r  $?  a    5  $  $?  0:  �E  r  $?  �x   5  �  $?  X:  �E  r  $?  �y   )z0  ]A  �<  �U  07  3  �:  @  @  ��   [	@  8�N   \$   ��<  �   $!,�  !-�  K  !:H<   �e  !=�   � !?�   "  !@�   �4  !A*>   �J  !B0>  �A  !O;  ;  6>   �A  !Q%;  0;  6>  <>   �A  !V@;  K;  6>  �    �
 !Y51  �:  c;  n;  B>  �:   �
 !]�R  �:  �;  �;  B>  �:   � !c?  �:  �;  �;  6>  �:  �   _ !m.   �;  �;  6>  �:  �:   �3  !q89  �:  �;  �;  B>   .E  !��3  <  <  6>  �:  0>   �(  !��(  3<  ><  6>  �:   ]_Tp H    �:  8ZD  88E  ^U  $A>  q<  �?  �    _9+  $N>  �?  �     �� \2*  7�<  `8.   a~  a�  �  �  ~  a�  �  8"�=  �{  "�   ]�  "�  \�  " �  �D  "!�  �3  ""�  U>  "#�  &�  "$�  �  "%�  �*  "&�   ڡ  "'H   $�U  "(H   %TL  ")H   &�I  "*H   'Q  "+H   (�C  ",H   )�J  "-H   *1  ".�  ,o(  "/H   0�U  "0H   1PL  "1H   2�I  "2H   3Q  "3H   4�C  "4H   5�J  "5H   6 W)%  "K�  >  �   �   bGT  "P>  �<  �  # �   aH   a�  �:  aH<  H<  �  az    �   �<  �      �  a�  a  a  cA   �>  d �  �  �>  �>  �    a�"  �"  E   a�"  �"  �>  �"  �  c�>  �>  d c?  ?  d ?  �>  a�"  �"  a�#  $?  a�&  �&  $'  e�   A?  f G?  g�5  6?  �&  �  r'  a�'  o?  ec?  ~?  c?   �?  e�?  �?  �?   a~'  �?  e?  �?  ?   �*  [  3  a[  a3  S3  @3  aw3  a@3  �4  >  hW<  @  iXF  $A�?  i\;  $A�   jk�T  $C>    R/  �4  lf-  8@  B@  mh  B@   $@  l�-  U@  _@  mh  B@   l�-  m@  w@  mh  B@   l�-  �@  �@  mh  B@   z/  �4  l[/  �@  �@  mh  �@   �@  l�/  �@  �@  mh  �@   l�/  �@  �@  mh  �@  n__n !�    @  lD	  A  A  mh  A   k>  l�	  $A  .A  mh  A   ]-  l�-  BA  UA  mh  UA  m#  [>   .A  l�'  hA  �A  mh  �A  m#  [>  m�!  �A   Q?  W?  h�  �A  jo__p ��    hq<  �A  iXF  $N�?  i\;  $N�    l�  �A  �A  mh  �A  p__a ��A   w>  N>  h�  B  n__c 	 B   �<  l�/  B  BB  mh  �@  n__c �z/  jq�&  ��/    h
  eB  rhR  	$eB  rmR  	$jB   �<  �<  h�4  �B  p__a K�"  p__b K�"   h�4  �B  p__a O�"  p__b O�"   h
5  �B  p__a ��#  p__b ��#   h$5  �B  p__a ��#  p__b ��#   aX5  a�#  h>5   C  p__a � C  p__b ��#   �B  �&  l$  9C  CC  mh  CC   %C  aw5  a�"  h]5  uC  p__a [uC  p__b [�"   NC  h|5  �C  p__a W�"   h�5  �C  p__a _�C  p__b _�"   NC  �#  l:$  �C  �C  mh  �C  r�6  v3  jq'U  x3    �C  l^$  D  D  mh  CC   l}$  D  =D  mh  �C  r�R  �3  jq'U  �3    �5  l�2  QD  gD  mh  gD  n__c aH    =D  l.  zD  �D  mh  UA   0  l�/  �D  �D  mh  �@  n__s ��D  n__n �3   l.  �D  �D  mh  UA  i�%  �$   lb*  �D  E  mh  �A  n__s 7�?  n__n 73  jq>*  9�5    l#0  )E  3E  mh  �@   l7.  AE  VE  mh  UA  i�%  �$   lV.  dE  nE  mh  B@   l'  |E  �E  mh  �E   0?  h�5  �E  !T  H   �E  r  i�3  �@  i�D  �@  jkZ*  ��<    s)  l�$  �E  F  mh  �C  r�%  B�#  jq'U  D�#    l�$  F  AF  mh  �C  r�%  S�#  r�?  S�#  jq'U  U�#    l�  OF  dF  mh  dF  iQ  ��   �?  lt.  wF  �F  mh  B@   lB0  �F  �F  mh  �@  iQ  �{0  i@  �$  i^F  ��$   h�5  G  !T  H   �E  r  i%  ,G  p__s -�  p__n -3  jk>*  2�5    $?  5  tA  v G  *G  mh  *G   
G  l>4  =G  GG  mh  GG   �?  l�  ZG  dG  mh  dG   �?  l�0  wG  �G  mh  �@  rj(  o0  r^F  �$   h6  �G  �$  	  i\C  ��G  i?)  ��G   �?  �?  a�5  h16  �G  �R  �2  p__f .=D   hO6  -H  !T  H   �E  r  r%  J-H  !T  H   �E  r   $?  l�.  @H  JH  mh  B@   hw6  �H  !T  H   �E  r  i%  9�H  p__n 93  jo__c >�  jk>*  A�     $?  h�6  �H  �E  r  r%  ��H  n__c �H   �E  r   $?  h'  �H  n__s 	�<   h�6  "I  �E  r  r%  "I  n__s �  �E  r   $?  a7  7  h�6  RI  �R  �0  p__f .-I   l�3  `I  uI  mh  uI  p__s �zI   �?  �?  l�0  �I  �I  mh  �I  n__s 	�0  r$  	�I  r�O  	1  n__v 	:    -I  ?  l1  �I  J  mh  �I  n__s #	�0  r$  #	J  r�O  #	1  n__v $	A    ?  lL1  ,J  fJ  mh  �I  n__s ��0  r$  �fJ  r�O  �1  n__v ��<   ?  l1  yJ  �J  mh  �I  n__s )	�0  r$  )	�J  r�O  )	1  n__v )	�    ?  l�1  �J   K  mh  �I  n__s -	�0  r$  -	 K  r�O  -	1  n__v .	%    ?  l�1  K  MK  mh  �I  n__s ^	�0  r$  ^	MK  r�O  ^	1  n__v ^	3    ?  l2  `K  �K  mh  �I  n__s b	�0  r$  b	�K  r�O  b	1  n__v c	,    ?  lK2  �K  �K  mh  �I  n__s w	�0  r$  w	�K  r�O  w	1  n__v x	�   ?  #   l,    L  L  mh  L  r4&  r�   �K  l0;  )L  <L  mh  <L  m#  [>   6>  lb  OL  bL  mh  bL  m#  [>   H>  l�:  uL  L  mh  <L   l1  �L  �L  mh  bL   l;  �L  �L  mh  <L  �L   <>  lG  �L  �L  mh  bL  p__a s�L   N>  l�  �L  �L  mh  A   u�  
M  M  mh  M  m#  [>   e>  �7  l7  6M  @M  mh  @M   "M  lm  SM  ]M  mh  A   l�  kM  ~M  mh  ~M  m#  [>   q>  l27  �M  �M  mh  @M   l^7  �M  �M  mh  @M   l}7  �M  �M  mh  @M   l�7  �M  �M  mh  @M   �4  l�4  �M  N  mh  N  r4&  :�   �M  l�$   N  *N  mh  CC   h�7  _N  !T  H   p__s p@3  i�+  p�  iR'  p�    l�2  mN  �N  mh  gD  n__c 3H    v_N  �T  ��   ��N  �N  wmN  � wvN  � vZA  bC  ��   ��N  �N  xhA     y4A  ��   ]xBA  !  z��  vZA  "Q  М+   �O  ZO  whA  � {ZA  ؜   ]PO  xhA  D  |4A  ؜�  ]xBA  c  }�  ~��N�   l�'  hO  �O  mh  �A  m#  [>  m�!  �O  i(  T]?   W?  vZO  �F  �%   ��O  �O  xhO  �  xzO  �  w�O  �5�/  ���  vZO  �  @��   ��O  aP  whO  � w�O  �{lD  L�=   U*P  xzD  �  }U� {4A  ��   ULP  wBA  s�}�� ���/  �Ɲc�   vZA  �I  Н   �|P  �P  whA  � wzA  � ��'  �   ��P  �P  �h  �A  � �$%  li?  ������� �   �(   �   ��P  Q  �h  �A  � �$%  u~?  � �2(   �   �#Q  @Q  �h  �A  � �$%  �?  � ��D  MN  @�V   �\Q  >R  w�D  � w�D  �w E  ��M�   �Q  �E    ��D  V�   9x�D  $  x�D  Z  x�D  z    �  x�D  �  x E  �  x�D  �  �  �E  ��D  m�   ;x�D  �  x�D  �  ��B  m�8  �1R  x�B  �  x�B     ~��6/      ��*  ���   �VR  FT  �h  �A  � �P  1T  ��*  �$  1  {E  ��   ۚR  x)E  ]   ��D  Ҟx  ��R  x�D  p  x�D  �  {�B  ڞ   ��R  x�B  p  x�B  �   ��6/   ��  �S  �WT  �3E  ��  �zS  xJE  �  xAE  �  {�B  �   �oS  xC  �  x	C     y�B  �   �x�B  �  x�B  /    ��w�   ���}�  �C�w�  �M���   �3E  !��  �T  xJE  C  xAE  o  {�B  )�   �T  xC  C  x	C  �  y�B  )�   �x�B  C  x�B  �    �H�w�   ��}�  �8���  �]���   �V�c�  �f�c�   \  % WT  8�  \T  aQT  ��*  p��   �zT  MV  �h  �A  ���  8V  ��&  �Z'  � {AF  ��   ��T  �XF  xOF  �   ��F  ��  ��T  ��F  ��F  ��F   x�F  V   �(  �U  �MV  �3E  ��H  ��U  xJE  i  xAE  �  {�B  ��   �vU  xC  i  x	C  �  y�B  ��   �x�B  i  x�B  �    ��w�   ���}�  �;�w�  �E���   �3E  �`  �V  xJE    xAE  -  {�B  �   �V  xC    x	C  V  y�B  �   �x�B    x�B  �    �@�w�   ��}�  �-���  �U���   �N�c�  �^�c�   \T  ��*  `��   �jV  �X  �h  �A  � �%  Z'  ���  �X  ��*  $  �  ���/   �V  �__p ^+  �H�iG  ���  ��G  w�G  �TxwG  �    ��D  Ǡ�  CW  x�D  �  x�D    {�B  Ϡ   �8W  x�B  �  x�B  #   �ܠ6/   ��  �W  ��X  �3E  ��  �W  xJE  7  xAE  c  {�B  ��   ��W  xC  7  x	C  �  y�B  ��   �x�B  7  x�B  �    ��w�   ��}�  �6�w�  �@���   �3E  �   fX  xJE  �  xAE  �  {�B  �   �[X  xC  �  x	C    y�B  �   �x�B  �  x�B  ;    �;�w�   ��}�  �(���  �P���   �I�c�  �Y�c�   \T  �+  `��   ��X  [  �h  �A  � �Q  "f'  ���J  "$  ��   �Z  ��*  $$  O  ���"   TY  �__p +^+  �T��F  ��8  ,��F  w�F  uw�F  V�W�x�F  �    ��D  ��P  ;�Y  x�D  �  x�D  �  {�B  ��   ��Y  x�B  �  x�B  �   �̡6/   �h  UZ  �[  �3E  ��  56Z  xJE  �  xAE    {�B  �   �+Z  xC  �  x	C  *  y�B  �   �x�B  �  x�B  Y    ���w�   �ߡ}�  �&�w�  �0���   �3E  ��  9�Z  xJE  m  xAE  �  {�B  	�   ��Z  xC  m  x	C  �  y�B  	�   �x�B  m  x�B  �    �+�w�   ���}�  ����  �@���   �9�c�  �I�c�   \T  l=+  [  2[  mh  �A  m#  [>  m�!  2[   W?  v[  +  P�%   �R[  v[  x[    x([    u�/  ��0  v[  �%  ���   ��[  �[  w[  � �lD  ��=   ��[  xzD  -  }�� �4A  �   ��[  wBA  s�}�� ��/  ��c�   l�&   \  \  mh  \  i%  /\   *?  $?  v�[  f)  �e   �>\  �\  w\  � w\  ���D  `��  9�\  ��D  ��D  {�B  `�   ��\  ��B  x�B  x   ~u�6/   �C�>R   l�&  �\  �\  mh  \  m#  [>   ��\  �  ��a   ��\  k]  w�\  � �E  ��	   �]  x)E  �   ��D  ã�  �`]  ��D  x�D  �  {�B  ˣ   �U]  ��B  x�B  �   �أ6/   ���X:   �*  �T  ��]  N`  �h  �A  � ��3  x]?  ���  C`  ��*  z$  �  ��$  {�&  �X��E  �  �	^  x�E  �  x�E    �  ��E  �W�0�g:    �0  �^  �N`  �3E  �P  ��^  xJE  r  xAE  �  {�B  ��   ��^  xC  r  x	C  �  y�B  ��   �x�B  r  x�B  �    ��w�   �Ф��  ��}�  �6�w�   �3E  �h  �*_  xJE  
   xAE  *   {�B  �   �_  xC  
   x	C  H   y�B  �   �x�B  
   x�B  j     �;�w�   ��D  ;��  �{_  ��D  x�D  ~   {�B  C�   �p_  ��B  x�B  �    �M�6/   ��\  P��  �`  x�\  �   �E  p�	   ��_  x)E  �    ��D  ���  �`  x�D  �   x�D  !  {�B  ��   �`  x�B  �   x�B  !   ���6/   �e�X:   }	�}٤��}�  �(���  �B���   ��c�   \T  �?*  P�i  �k`  �c  �h  �A  � �__c �B'  ���  �c  ��$  ��&  �X��  	c  ��*  �$  /!  �  xa  k>*  �c+  |B  ~�0  �x'B  s!  xB  �!  �~�   *a  �4B  �!  ��@  ��   ���@  x�@  �!    � �   x'B  �!  xB  "  � �   �4B  ��A  �H  �w�A  �C�        ��D  �`  ��a  x�D  ("  x�D  <"  {�B  %�   ��a  x�B  ("  x�B  O"   �2�6/   �x  wb  ��c  �3E  P��  �Xb  xJE  c"  xAE  �"  {�B  V�   �Mb  xC  c"  x	C  �"  y�B  V�   �x�B  c"  x�B  �"    �e�w�   �N�}�  �j���  ���w�   �3E  ���  ��b  �JE  xAE  �"  {�B  ��   ��b  �C  x	C  #  y�B  ��   ���B  x�B  /#    ���w�   ���}�  �����  �����   ��\  ���  ��c  x�\  C#  �E  ��	   �Ec  x)E  #   ��D  ӥ�  ��c  x�D  �#  x�D  �#  {�B  ۥ   ��c  x�B  �#  x�B  �#   ��6/   ���X:   }i�}s� �{�c�   \T  ��*  ��B  ��c  g  �h  �A  � �__s ��  ��__n �3  ���  g  ��$  ��&  �X{�D  �7   �e  x E  �#  x�D  <$  x�D  h$  ��   �d  �E  �$  ��D  �   9x�D  �$  x�D  %  x�D  J%    ���   x�D  ]%  x E  q%  x�D  �%  ���   �E  ��D  �   ;x�D  �%  x�D  �%  {�B  	�   �e  x�B  �%  x�B  �%   ��6/      �8  �e  �g  �3E  ��P  Ǩe  xJE  �%  xAE  �%  {�B  ��   ��e  xC  �%  x	C  &  y�B  ��   �x�B  �%  x�B  2&    ���w�   ���}�  �ڧw�  �ߧ��   �3E  ��h  �@f  xJE  F&  xAE  f&  {�B  ��   �5f  xC  F&  x	C  �&  y�B  ��   �x�B  F&  x�B  �&    ���w�   ��\  ��  ��f  x�\  �&  �E  9�	   �|f  x)E  �&   ��D  c��  ��f  x�D  	'  x�D  '  {�B  k�   ��f  x�B  	'  x�B  0'   �x�6/   �.�X:   }٦���}�  �̧��  }�� ���   ��c�   \T  vnE  �3  �   �3g  <g  w|E  �  l�.  Jg  `g  mh  B@  n__c �H    �8   �s   �ch  !T  H   �E  r  �%  4ch  � �<g  +��  50h  �Sg  
xJg  D'  ��G  2��  ��g  x�G  �'  ����:   �CD  6��  �xZD  �'  xQD  �'  �`�.   xZD  �'  xQD  �'  �i��2     ��G  J� 	  5Xh  xH  �'  ~X�>R   �J�S`   $?  �78  ��   ��h  !T  H   �E  r  �%  @�h  � ���S`   $?  ��G  m   ��   ��h  wH  � Ũ>R  �� �   l�.  �h  i  mh  UA  r�R  ��.  jq'U  ��.    �c8  Шz   �>j  !T  H   �E  r  �%  
�>j  
(  �__f 
�3  @(  |�h  ި	  
�w�h  �x�h  �(  �	  �i  �(  �2H  ި8	  �x@H  �(  �<g   �`	  p�Sg   xJg  �(  ��G  �x	  ��i  x�G  �(  �J��:   �CD  ��	  �xZD  	)  xQD  )  � �%   xZD  <)  xQD  Q)  �)��2         $?  ��8  P�   �k  !T  H   �E  r  �%  
mk  � �__f 
m�,  d)  y�E  ]�   
ow�E  �w�E  R�]�   ��E  �)  �TC  ]�   EwiC  �w^C  r�y�B  ]�   \w�B  �x�B  �)       $?  ��8  p�   ��k  !T  H   �E  r  �%  
O�k  � �__f 
O�,  �|F  y��	  
Qx&F  �)  �F   wF  Q��	  �3F  �)  �zC  y��	  V�k  x�C  �)   ��C  ��   Vx�C  �)  w�C  q�yoB  ��   `x�B  �)  xyB  �)       $?  ��8  ��G   �m  !T  H   �E  r  �%  
�m  �)  �__f 
�-  
*  yF  ��   
�x&F  4*  �F  xF  I*  ���   �3F  r*  ��C  ��   V�l  x�C  �*  x�C  �*  yoB  ��   `x�B  �*  xyB  r*    �TC  ��   WxiC  �*  x^C  �*  y�B  ��   \x�B  �*  x�B  �*       $?  �#9  �   �~m  !T  H   �E  r  �%  
�~m  � �__f 
�+-  +  |�C  ��	  
�x�C  /+  w�C  ���	  ��C  ^+     $?  �S9   �   ��m  !T  H   �E  r  �%  
��m  � �__f 
�D-  }+  |D  ��	  
�xD  �+  w"D  ���	  �/D  �+     $?  ��9   �   ��v  !T  H   �E  r  �%  L�v  � �__s M�  ��__n M3  ��
  �v  ��$  R�&  �X�0
  �t  o__w W�5  �P
  �s  ��-  Z`>  �+  {oB  U�   [�n  x�B  �,  xyB  �,   {�F  #�1   `�o  x�F  	-  ��F  x�F  -  �#�   -o  ��F  \-  y�D  #�   2x�D  o-  ��D  x�D  �-    �:�   ��F  ��F  x�F  �-  �:�   ��F  |�D  <�p
  4x�D  �-  x�D  �-  {�B  D�   ��o  x�B  �-  x�B  �-   �Q�6/      �JH  u��
  b�q  xqH  �-  xfH  .  ��
  Dq  �}H  C.  �2H  u��
  >�p  x@H  W.  �<g  ��  pxSg  �.  xJg  �.  ��G  ��@  �Tp  x�G  H/  �{��:   �CD  ��`  �xZD  �/  xQD  �/  ��  xZD  0  xQD  60  �+��2      ��  ��H  |B  ���  Ax'B  V0  xB  v0  ��  q  x'B  �0  xB  �0  ��  �4B  ��A  ��   �x�A  �0     ��  �4B  �0  ��@  ��   ���@  x�@  �0       �֫
   �qH  xfH  �0  �֫
   �}H  �֫
   ��H      |JH  ��  ^xqH  1  xfH  �1  �   s  �}H  �1  �2H  �H  >hr  x@H  �1  �<g  �p  pxSg  j2  xJg  �2  ��G  ���  �r  x�G  �2  �v��:   �CD  ���  �xZD  33  xQD  b3  ��  xZD  �3  xQD  �3  �Y��2      ��  ��H  |B  ���  Ax'B  �3  xB  �3  �  �r  x'B  4  xB  %4  �  �4B  ��A  ��   �x�A  84     �(  �4B  P4  ��@  �   ���@  x�@  c4       �F�*   �qH  xfH  w4  �F�*   �}H  �F�*   ��H  |�D  H�@  Dx�D  �4  x�D  �4  {�B  P�   ��s  x�B  �4  x�B  �4   �]�6/        {�F  ӪP   e�t  x�F  �4  x�F  �4  x�F  �4  �X  t  ��F   5  y�D  Ӫ   2x�D  5  x�D  '5  x�D  ;5    �p  ��F  ��F  x�F  N5  �p  ��F  y�D  ��/   4x�D  l5  x�D  �5  {�B  ��   �{t  x�B  l5  x�B  �5   ��6/      yD  ��   fxD  �5  x"D  �5  ���   �/D  �5     ��  iu  ��v  �3E  ���  jJu  xJE  �5  xAE  6  {�B  ��   �?u  xC  �5  x	C  +6  y�B  ��   �x�B  �5  x�B  Z6    �ŭw�   ���}�  ���w�  �����   �3E  Э�  n�u  xJE  n6  xAE  �6  {�B  ح   ��u  xC  n6  x	C  �6  y�B  ح   �x�B  n6  x�B  �6    ��w�   ��\  ���  p�v  x�\  �6  �E  ��	   �v  x)E  7   ��D  s��  �vv  x�D  17  x�D  E7  {�B  {�   �kv  x�B  17  x�B  X7   ���6/   ���X:   }6��έ}�  ����  }�����   ��c�   $?  \T  ��H  $   �   ��v  w�H  � w�H  ��;� n   ��9  @�   �]w  �E  r  �%  �]w  � �__c �Z   ���H  K�   �x�H  l7  w�H  � �[� n    $?  ��9  `�   ��w  �E  r  �%  ��w  � �__c �a   ���H  k�   �x�H  �7  w�H  � �{� n    $?  ��H  �/  ��R   ��x  w I  � wI  ���H  ��   #x  x�H  �7  �����   ���   �x  �I   x I  �7  ��D  ��  ��D  x�D  �7  {�B  ��   ��x  ��B  x�B  8   �Ǯ6/    ��� n   �x  Z   �:  �R   ��y  �E  r  �%  $�y  � �__s $�x  ���H  �   %xI  &8  x I  \8  ��H  �   1y  x�H  �8  �����   ��   �y  �I   x I  �8  ��D  �8  ��D  x�D  �8  {�B  �   ��y  ��B  x�B  �8   �'�6/    �� n    $?  �y  a   �0:  @�R   ��z  �E  r  �%  �z  � �__s �y  ���H  M�P   xI  �8  x I  +9  ��H  Q�   Ez  x�H  `9  �Z���   �p�   �z  �I   x I  9  ��D  r�h  ��D  x�D  �9  {�B  z�   ��z  ��B  x�B  �9   ���6/    �e� n    $?  �h+  ��  ��z  �~  ]T  :   �h  �A  � �__v @:   ���  �~  ��$  B�&  �X��  ~  ��*  E$  �9  ��  �|  ��#  H�~  :  �3I  ̯�  Hw{  xFI  H:  �'��:   �2H  ԯ  I-|  x@H  �:  �<g  p�0  pxSg  �:  xJg  �:  ��G  s�P  ��{  x�G  ;  �.��:   �CD  ~�p  �xZD  m;  xQD  �;  ��B   xZD  �;  xQD  �;  ���2      {RI  �   IP|  xiI  �;  �`I   yI  �   Ix�I  <  ��I  x�I  v<  x�I  �<  x�I  �<    ��D  ��  T�|  x�D  �<  x�D  �<  {�B  �   ��|  x�B  �<  x�B  �<   �'�6/   ��  �}  ��~  �3E  B��  Nk}  xJE  �<  xAE  =  {�B  H�   �`}  xC  �<  x	C  -=  y�B  H�   �x�B  �<  x�B  O=    �W�w�   �@�}�  �\���  �y�w�   �3E  ���  R�}  �JE  wAE  W{�B  ��   ��}  �C  w	C  w�y�B  ��   ���B  x�B  c=    ���w�   ���}�  �����  �����   ��\  *��  V�~  x�\  w=  �E  J�	   �V~  x)E  �=   ��D  ��  ��~  x�D  �=  x�D  �=  {�B  ��   ��~  x�B  �=  x�B  �=   �Ȱ6/   �?�X:   }��}h� �p�c�   �~  a�+  \T  �U(  ��   ��~  0  �h  �A  � �__n �:   ����z  �� � ���  ��(  ��@   �H  �  �h  �A  >  �__n \o   +>  �ȱ8   k-  `%  {oB  ͱ   `�  ��B  JxyB  K>   ~��z  ~ ��z    �)   �   ��  �  �h  �A  � �__n j�   �� �   k-  n%  ��z  �� � ���   ��+  �  �;�  $�  ]T  A   �h  �A  � �__v @A   ��   �  ��$  B�&  �X�H  o�  ��*  E$  >  �p  ��  ��#  H$�  �>  �3I  <��  H̀  xFI  ?  ����:   �2H  D��  I��  x@H  B?  �<g  ��  pxSg  v?  xJg  �?  ��G  ��  �5�  x�G  �?  ����:   �CD  �  �xZD  (@  xQD  J@  �P�B   xZD  �@  xQD  �@  �[��2      {RI  Z�   I��  xiI  �@  �`I   y�I  ^�   IxJ  �@  � J  x�I  1A  x�I  DA  x�I  \A    ��D  ��(  T7�  x�D  oA  x�D  �A  {�B  ��   �,�  x�B  oA  x�B  �A   ���6/   �@  ߂  �)�  �3E  ��X  N��  xJE  �A  xAE  �A  {�B  ��   ���  xC  �A  x	C  �A  y�B  ��   �x�B  �A  x�B  
B    �ǳw�   ���}�  �̳��  ��w�   �3E  ��p  RP�  �JE  wAE  W{�B  ��   �E�  �C  w	C  w�y�B  ��   ���B  x�B  B    ��w�   ��}�  ����  ����   ��\  ���  V�  x�\  2B  �E  ��	   ���  x)E  nB   ��D  #��  ��  x�D  �B  x�D  �B  {�B  +�   ���  x�B  �B  x�B  �B   �8�6/   ���X:   }&�}س ��c�   �~  \T  �x(   �   �F�  �  �h  �A  � �__n �A   �%��  �� � ���  ��(  0�   ���  Ȅ  �h  �A  � �__n �h   �B  >��  �� �   �')  @�   ���  �  �h  �A  � �__n �v   �E��  �� � ���  ��+  P�  �:�  #�  ]T  �<  �h  �A  � �__v @�<  ���  �  ��$  B�&  �X��  n�  ��*  E$  �B  �  ݆  ��#  H#�  +C  �3I  ��(  H˅  xFI  _C  ���:   �2H  ��@  I��  x@H  �C  �<g  0�h  pxSg  �C  xJg  �C  ��G  3��  �4�  x�G  D  ���:   �CD  >��  �xZD  nD  xQD  �D  ���B   xZD  �D  xQD  �D  ����2      �J  ���  I��  xYJ  �D  �MJ  xAJ  E  �5J  x,J  #E   yRI  ��   IxiI  6E  �`I    ��D  ״�  T4�  x�D  IE  x�D  ]E  {�B  ߴ   �)�  x�B  IE  x�B  pE   ��6/   ��  ܇  �(�  �3E  �  N��  xJE  �E  xAE  �E  {�B  �   ���  xC  �E  x	C  �E  y�B  �   �x�B  �E  x�B  �E    ��w�   � �}�  ����  �9�w�   �3E  D�   RO�  �JE  xAE  F  {�B  L�   �D�  �C  x	C  .F  y�B  L�   ���B  x�B  PF    �e�w�   �B�}�  �[���  �l���   ��\  �@  V�  x�\  dF  �E  �	   ���  x)E  �F   ��D  s�X  ��  x�D  �F  x�D  �F  {�B  {�   ���  x�B  �F  x�B  �F   ���6/   ��X:   }l�}(� �0�c�   �~  \T  ��(  p�   �E�  v�  �h  �A  � �__n ��<  �F  ~��  �� �   ��+  ��  ���  ��  ]T  �   �h  �A  � �__v @�   ��p  u�  ��$  B�&  �X��  ˌ  ��*  E$  G  ��  <�  ��#  H��  ]G  �3I  ���  H(�  xFI  �G  ���:   �2H  ���  Iފ  x@H  �G  �<g  `�   pxSg  H  xJg  3H  ��G  c�@  ���  x�G  \H  ���:   �CD  n�`  �xZD  �H  xQD  �H  �зB   xZD  I  xQD  0I  �۷�2      {RI  ֶ   I�  xiI  DI  �`I   ykJ  ڶ   Ix�J  WI  ��J  x�J  kI  x�J  ~I  xyJ  �I    ��D  ��x  T��  x�D  �I  x�D  �I  {�B  �   ���  x�B  �I  x�B  �I   ��6/   ��  ;�  ���  �3E  2��  N�  xJE  �I  xAE  J  {�B  8�   ��  xC  �I  x	C  "J  y�B  8�   �x�B  �I  x�B  DJ    �G�w�   �0�}�  �L���  �i�w�   �3E  t��  R��  �JE  wAE  W{�B  |�   ���  �C  w	C  w�y�B  |�   ���B  x�B  XJ    ���w�   �r�}�  �����  �����   ��\  ��  Vj�  x�\  lJ  �E  6�	   ��  x)E  �J   ��D  ���  �_�  x�D  �J  x�D  �J  {�B  ��   �T�  x�B  �J  x�B  �J   ���6/   �+�X:   }��}X� �`�c�   �~  \T  �J)  ��   ���  ݍ  �h  �A  � �__n ɚ   ���v�  �� � ����%  �,  ��  ���  �  ]T  %   �h  �A  � �__v @%   ��  ܑ  ��$  B�&  �X�8  2�  ��*  E$  �J  �`  ��  ��#  H�  FK  �3I  ��  H��  xFI  zK  �G��:   �2H  ��  IE�  x@H  �K  �<g  ���  pxSg  �K  xJg  L  ��G  ���  ���  x�G  EL  �N��:   �CD  ��   �xZD  �L  xQD  �L  � �B   xZD  M  xQD  M  ���2      {RI  �   Ih�  xiI  -M  �`I   y�J  
�   Ix�J  @M  ��J  x�J  TM  x�J  gM  x�J  M    ��D  .�  T��  x�D  �M  x�D  �M  {�B  6�   ��  x�B  �M  x�B  �M   �C�6/   �0  ��  ��  �3E  b�H  N��  xJE  �M  xAE  �M  {�B  h�   �x�  xC  �M  x	C  N  y�B  h�   �x�B  �M  x�B  -N    �w�w�   �`�}�  �|���  ���w�   �3E  ��`  R�  �JE  wAE  W{�B  ��   ��  �C  w	C  w�y�B  ��   ���B  x�B  AN    �źw�   ���}�  �����  �̺��   ��\  F��  Vё  x�\  UN  �E  f�	   �n�  x)E  �N   ��D  ӹ�  �Ƒ  x�D  �N  x�D  �N  {�B  ۹   ���  x�B  �N  x�B  �N   ��6/   �[�X:   }Ҹ}�� ���c�   �~  \T  �m)  к   �	�  D�  �h  �A  � �__n �%   �պݍ  �� � ����%  �I,  �  �e�  N�  ]T  3   �h  �A  � �__v @3   ���  C�  ��$  B�&  �X��  ��  ��*  E$  �N  �  
�  ��#  HN�  /O  �3I  �(  H��  xFI  cO  �g��:   �2H  �@  I��  x@H  �O  �<g  ��h  pxSg  �O  xJg  P  ��G  ���  �_�  x�G  .P  �n��:   �CD  ���  �xZD  �P  xQD  �P  � �B   xZD  �P  xQD  Q  �+��2      {RI  0�   Iϓ  xiI  Q  �`I   yK  4�   Ix@K  )Q  �4K  x(K  =Q  xK  PQ  xK  hQ    ��D  X��  Ta�  x�D  {Q  x�D  �Q  {�B  `�   �V�  x�B  {Q  x�B  �Q   �m�6/   ��  	�  �S�  �3E  ���  N�  xJE  �Q  xAE  �Q  {�B  ��   �ߔ  xC  �Q  x	C  �Q  y�B  ��   �x�B  �Q  x�B  R    ���w�   ���}�  �����  ���w�   �3E  ļ  Rz�  �JE  wAE  W{�B  ̼   �o�  �C  w	C  w�y�B  ̼   ���B  x�B  *R    ��w�   �¼}�  �ۼ��  ����   ��\  p�(  V8�  x�\  >R  �E  ��	   �Օ  x)E  zR   ��D  �@  �-�  x�D  �R  x�D  �R  {�B  ��   �"�  x�B  �R  x�B  �R   ��6/   ���X:   }��}�� ���c�   �~  \T  ��)  �   �p�  ��  �h  �A  � �__f �3   ���D�  �� � ����3  ��)   �   �Ö  �  �h  �A  � �__f ��<  ���D�   �u,   �  ��  ��  ]T  ,   �h  �A  � �__v @,   ��X  �  ��$  B�&  �X��  ?�  ��*  E$  �R  ��  ��  ��#  H��  S  �3I  L��  H��  xFI  LS  ����:   �2H  T��  IR�  x@H  �S  �<g  �  pxSg  �S  xJg  �S  ��G  �(  ��  x�G  T  ����:   �CD  ��H  �xZD  qT  xQD  �T  �`�B   xZD  �T  xQD  �T  �k��2      {RI  j�   Iu�  xiI  �T  �`I   yRK  n�"   Ix�K  U  ��K  xuK  &U  xiK  9U  x`K  QU    ��D  ��`  T�  x�D  dU  x�D  xU  {�B  ��   ���  x�B  dU  x�B  �U   ���6/   �x  ��  ���  �3E  ¾�  N��  xJE  �U  xAE  �U  {�B  Ⱦ   ���  xC  �U  x	C  �U  y�B  Ⱦ   �x�B  �U  x�B  �U    �׾w�   ���}�  �ܾ��  ���w�   �3E  ��  R �  �JE  wAE  W{�B  �   ��  �C  w	C  w�y�B  �   ���B  x�B  V    �%�w�   ��}�  ����  �,���   ��\  ���  Vޚ  x�\  'V  �E  н	   �{�  x)E  cV   ��D  3��  �Ӛ  x�D  vV  x�D  �V  {�B  ;�   �Ț  x�B  vV  x�B  �V   �H�6/   �ŽX:   }6�}� ��c�   �~  \T  ��)  0�   ��  Q�  �h  �A  � �__f �,   �5��  �� � ����,  ��,  @�  �r�  [�  ]T  �  �h  �A  � �__v @�  ���  P�  ��$  B�&  �X�   ��  ��*  E$  �V  �H  �  ��#  H[�  W  �3I  l�h  H�  xFI  5W  ����:   �2H  t��  I��  x@H  tW  �<g  ��  pxSg  �W  xJg  �W  ��G  ��  �l�  x�G   X  ����:   �CD  ��  �xZD  ZX  xQD  |X  ���B   xZD  �X  xQD  �X  ����2      {RI  ��   Iܜ  xiI  �X  �`I   y�K  ��   Ix�K  �X  ��K  x�K  cY  x�K  vY  x�K  �Y    ��D  ��   Tn�  x�D  �Y  x�D  �Y  {�B  ��   �c�  x�B  �Y  x�B  �Y   �ǿ6/   �  �  �`�  �3E  ��0  N��  xJE  �Y  xAE  �Y  {�B  ��   ��  xC  �Y  x	C  Z  y�B  ��   �x�B  �Y  x�B  <Z    ���w�   ���}�  �����  ��w�   �3E  $�H  R��  �JE  wAE  W{�B  ,�   �|�  �C  w	C  w�y�B  ,�   ���B  x�B  PZ    �E�w�   �"�}�  �;���  �L���   ��\  ʿh  VE�  x�\  dZ  �E  �	   ��  x)E  �Z   ��D  S��  �:�  x�D  �Z  x�D  �Z  {�B  [�   �/�  x�B  �Z  x�B  �Z   �h�6/   �߿X:   }V�}� ��c�   �~  \T  ��)  P�   �}�  ��  �h  �A  � �__p ��  �U�Q�  �� � ���  �U  =ß   �   ��   >ß  �B  ?ß  ��  E�   �   �B   F�  �C  G�  �e  H�  �8  I�  ��  J�  �

  XB�   �   ��  YB�  ��
  ZB�  ��   `n�  �   ��  f��   �   ��  g��  ��  h��  ��  n��   �   ��	  o��  ��  p��  �H  vؠ   �   �`  wؠ  �w  xؠ  �   yؠ  �~  �   �   �   ��  ��  ��  �  ��  ��   ��  ��  ��  ��	  ��  ��  �q�   �   �  �q�  �  �q�  ��  �q�  ��  ���     ��  ���  ��  ���  ��  ���  �m  ��     �	  ��  �2	  ��  ��  ��  �9  ��  �[  �)�     �J  �)�  ��  �)�  �7  �)�  ��  �b�   %  �I	  �b�  �$	  �b�  ��   ���   0  �N  ���  �p  ���   ;  ��  ���  �:  ���  ��  ­�  �d   í�  ��  ��   F  �  ��  ��  ��  ��	  ��   Q  ��  ��  �  �>�   \  ��  �>�  ��  �>�  ��  �>�  �+  �w�   g  ��  �w�  ��   �w�  �  飣   r  ��
  ꣣  ��  룣  �  �ϣ   }  �   �ϣ  �F  �ϣ  ��  ���   �  ��  ���  ��  ���  �D  O'�   �  ��  P'�  �1  Q'�  ��  WS�   �  �^  XS�  ��  3r�   �  ��  4r�  ��   8��   �  ��  9��  �l	  =��  �  �N  >��  �^  ?��  �L  @��  �a  D�  �  �B  E�  ��	  F�  �  G�  �  H�  �y  I�  ��   <�   �  ��  !<�  �  &�1  c�  �   �>  Y  w�  �   ��  ��  �  ��  �   ��  a�<  �O2  Y2  A   �    '>   �  �]  [  �V  �      +&  std # �   %  0
@?)  �=  �  �b  �%  Fe  �N%  �3  �=  z   J)  P)   	J   
eq �<-  V)  �   P)  P)   
lt ��1  V)  �   P)  P)   ��  eF  N%  �   ])  ])  �   �K  �9  �  �   ])   �(  
!  ])    ])  �  P)   1  �A  c)  ?  c)  ])  �   �5  �'  c)  c  c)  ])  �   �3  �A  c)  �  c)  �  J    +  :  J   �  i)   	U   �C   �P  U   �  P)   �B  $6  V)  �  i)  i)   eof (�:  U   ?  ,N0  U   i)    E  �  9Q  pz  G0  sz   �T  t?)  %  {E  K  �-   %  �[  f  �-  z   �:  �b;  z  ~  �  �-   �T  �4>  �  �  �-  ?)   �T  �QM  ?)  �  �  �-   �F  ��?  �-  �  �  �-  z    I  �O  �-  �    �-  z   (*  �	H      *  �-  z   �O  �eT    B  M  �-  z   �O  ́?  z  e  p  �-  �-   �$  ?)   �:  Z\%  _� �2%  �?  �U%  K  	\  �    �e  	_�  �4  	co)  �J  	du)  ��  	q�  �  �)   ��  	s�    �)  �)   W  	y  �)  N%    	�  5�)  6�*  7�*  �J  p�  �B  ~  �   %  �&   �B  m  +  �&  �)    �e  y�  [V  �  	~  �G  !A   <  x�  �4  {�  �J  |�  �J  {"  `S  ��"  ~J  ��  �J  ��  �%  �.  �K  �~   I  �~  :!  ��*   %H  ��  �   �3  2�  �G  7)  t3  B2+  �'  ��O   +  V  ��N  V)  �  �  =+   3  �o+  V)  �  �  =+    �P  ��O  �  �  +    �M  ��P  �  �  +    �,  �-  �  �  +  ~   �+  ��R  �&      +   3  �   �&  .  >  +  �)  �)   �/  !�B  +  b  ~  ~  �)    �O  �|6  u  �  +  �)   !(  ��6  �  �  +  �)   "�   �-  �&  �  �  +   #�1  o�*  �&  �  +  �)  ~    "�A  $n%  �&  �     +   "�A  (�I  �&    #  +  �&   ""A  ,�%  +  ;  A  +   "�1  2E)  �  Y  _  +   "�/  6;&  �  w  }  +   !�>  :�>  �  �  +   "S  A:2  ~  �  �  +  ~  )   !�#  K�(  �  �  +  ~  ~  )   "9  S>$  ~       +  ~  ~   "-U  [�7  V)  (  3  +  )   $�5  d�-  S  �&  )  ~   $	1  m�P  s  �&  )  ~   $�3  v\-  �  �&  ~  �%   $nU  ��-  �  �&  �  �   $nU  �nG  �  �&  �  �   $nU  ��   �  �&  �&  �&   $nU  �IP  	  �&  )  )   �J  �rR  N%  2	  ~  ~   !�=  ��H  F	  [	  +  ~  ~  ~   !V  �)  o	  u	  +   %�'  �D*   +  &�0  ��	  �	  +   '�0  ��	  �	  +  �)   �0  ��	  �	  +  &+   �0  ��	  �	  +  &+  ~  ~   �0  �
  !
  +  &+  ~  ~  �)   �0  �1
  F
  +  )  ~  �)   �0  �V
  f
  +  )  �)   �0  �v
  �
  +  ~  �%  �)   &�0  "�
  �
  +  N%   (�  *,Q  ,+  �
  �
  +  &+   (�  2�G  ,+  �
  �
  +  )   (�  =�%  ,+      +  �%   (S� f�&  �  ,  2  +   (S� q�>  �  K  Q  +   )end y<  �  j  p  +   )end �6;  �  �  �  +   (I ��$  �  �  �  +   (I ��7  �  �  �  +   (��  �lC  �  �  �  +   (��  �CM  �      +   (r ��R  ~  $  *  +   (�K  �r5  ~  C  I  +   (�3  �j=  ~  b  h  +   *�� �  }  �  +  ~  �%   *�� ��F  �  �  +  ~   (I  v  ~  �  �  +   *�E  �|U  �  �  +  ~   *�1  -�      +   (�� 5�?  V)     &  +   (�:  D�6  �  ?  J  +  ~   (�:  UW  �  c  n  +  ~   )at k
/  �  �  �  +  ~   )at ��7  �  �  �  +  ~   (�F  ��/  ,+  �  �  +  &+   (�F  �k:  ,+  �  �  +  )   (�F  ��H  ,+       +  �%   (@  DA:  ,+  9  D  +  &+   (@  U�1  ,+  ]  r  +  &+  ~  ~   (@  )�D  ,+  �  �  +  )  ~   (@  ��*  ,+  �  �  +  )   (@  �6  ,+  �  �  +  ~  �%   *�G  -aN  �    +  �%   �3  �b*  ,+     +  +  &+   (�3  ^ 2  ,+  D  Y  +  &+  ~  ~   (�3  �=  ,+  r  �  +  )  ~   (�3  z�T  ,+  �  �  +  )   (�3  � @  ,+  �  �  +  ~  �%   *� ��E  �  �  +  �  ~  �%   (� �\+  ,+    "  +  ~  &+   (� �u>  ,+  ;  U  +  ~  &+  ~  ~   (� g|=  ,+  n  �  +  ~  )  ~   (� "�@  ,+  �  �  +  ~  )   (� 9k<  ,+  �  �  +  ~  ~  �%   (� K�'  �  �    +  �  �%   (bL  d�R  ,+    ,  +  ~  ~   (bL  t�2  �  E  P  +  �   (bL  �L&  �  i  y  +  �  �   (�%  �9F  ,+  �  �  +  ~  ~  &+   (�%  �|<  ,+  �  �  +  ~  ~  &+  ~  ~   (�%  ��T  ,+  �    +  ~  ~  )  ~   (�%  ��A  ,+  +  @  +  ~  ~  )   (�%  b>  ,+  Y  s  +  ~  ~  ~  �%   (�%  3%  ,+  �  �  +  �  �  &+   (�%  'V7  ,+  �  �  +  �  �  )  ~   (�%  <�+  ,+  �    +  �  �  )   (�%  Q'S  ,+    5  +  �  �  ~  �%   (�%  vj.  ,+  N  h  +  �  �  �&  �&   (�%  ��9  ,+  �  �  +  �  �  )  )   (�%  �C  ,+  �  �  +  �  �  �  �   (�%  �>/  ,+  �    +  �  �  �  �   "�?  ��&  ,+    3  +  ~  ~  ~  �%   "�1  �O  ,+  K  e  +  ~  ~  )  ~   ,)  �z-  �&  �  ~  �%  �)   ++E  �3J  �&  �  ~  �%  �)   (�5  ��)  ~  �  �  +  �&  ~  ~   *n	 @D  �  �  +  ,+   (W�  �6  )      +   (�A  %�A  )  2  8  +   (��  ,Z5  �  Q  W  +   (�(  �;  ~  p  �  +  )  ~  ~   (�(  I�%  ~  �  �  +  &+  ~   (�(  X�5  ~  �  �  +  )  ~   (�(  �^   ~  �     +  �%  ~   (�(  v�S  ~    )  +  &+  ~   (�(  	K  ~  B  W  +  )  ~  ~   (�(  �o?  ~  p  �  +  )  ~   (�(  J5  ~  �  �  +  �%  ~   (NW  ��Q  ~  �  �  +  &+  ~   (NW  /�I  ~  �     +  )  ~  ~   (NW  ��,  ~    )  +  )  ~   (NW  ��;  ~  B  R  +  �%  ~   (�S  ��I  ~  k  {  +  &+  ~   (�S  >T?  ~  �  �  +  )  ~  ~   (�S  05  ~  �  �  +  )  ~   (�S  $S:  ~  �  �  +  �%  ~   (�>  2hL  ~    $  +  &+  ~   (�>  SUB  ~  =  R  +  )  ~  ~   (�>  Q�2  ~  k  {  +  )  ~   (�>  _�K  ~  �  �  +  �%  ~   (�4  qT  ~  �  �  +  &+  ~   (�4  j�K  ~  �  �  +  )  ~  ~   (�4  ��5  ~    $  +  )  ~   (�4  N.  ~  =  M  +  �%  ~   (U+  �)  5  f  v  +  ~  ~   (��  �!1  N%  �  �  +  &+   (��  ��T  N%  �  �  +  ~  ~  &+   (��  ��O  N%  �     +  ~  ~  &+  ~  ~   (��  �;.  N%    $  +  )   (��  ��B  N%  =  R  +  ~  ~  )   (��  ��,  N%  k  �  +  ~  ~  )  ~   	.  !T  �%  ,�E  >   ,�F  �   -�&  -�7  	5  .W  3D  /�4  /�$  /q-  /c=  /o'  /�5   /�%  � /�8  �/X)  �/�%  �/�  �/aO  �/Y=  � /P  �� /�C  ��/wS  �/�O  � /�?  �/�5  �� .
$ g}  /)W  /�   /�U  /�A  /�8  /�P   /EH  �� .�4  ��  /O   /�7  /(  /�Q  /G  �� .��  ��  /�R   /�-  /�1  /lO  �� 0b4 �  1�N  ��  1�9  iD  �P  ��  2�4    	�  3dec   2t-    3hex   2r'    2<    3oct   @2�   �4[)     4�%  "   4�  &   4dO  )   4\=  ,   4�P  /    4�C  3   @2zS  6  �2�O  9  J4�?  <  1�  J}  2�7  N$  		  2(  Q$  2�Q  V$  2O  Y$   3in w`  	�  3out z`  3beg ��   	�  3cur ��   0�8  �  !T  �%  ,�E  >    0�Y  �  !T  �%  ,�E  >    0�M     5Z  ��  �  �  6.  N%   &�B �    6.   !T  �%  ,�E  >    0�+  �  (��  a�)  M  B  M  �.  �%   1�b  ��%  6KC  3�T  M     {  �  �.  �%   7+3  ��3  �  �.    bH'  cO+  eZ+  fr+  g�+  h�+  i�+  j�+  k�+  l�+  m,  q9,  r^,  t},  u�,  v�,  x�,  y�,  |�,  ~-  �"-  �7-  �Q-  �c-  �y-  ��-  ��-  ��-  	  �^  -H'  �>  b�  	   8N  .?0  �  �R     �.   �\  �
K[  C+  �  !T  �%  �E  >   �F  �  C+  &+   0�E  %   (��  ��$     �     �6  �%   �b  K�%  !T  �%  ,�E  >    	�  t\  �
�[  I+  d   !T  �%  �E  >   �F  �  I+  ,+   +�V  L�L  C+  �   !T  �%  �E  >   C+  )  q   9	@  8�N  t\  �Z  I+  I+  ,+  �%    :$   E%  �  $,�  -�  K  :v"  �e  =�  � ?�&  "  @)  �4  Ao)  �J  Bu)  �A  O=!  C!  {)   �A  QS!  ^!  {)  �)   �A  Vn!  y!  {)  N%   �
 Y51  �   �!  �!  �)  !   �
 ]�R  	!  �!  �!  �)  !!   � c?  �   �!  �!  {)  �   �(   _ m.   �!  "  {)  �   �    �3  q89  �   #"  )"  �)   .E  ��3  ="  M"  {)  �   u)   �(  ��(  a"  l"  {)  �    ;_Tp �%   	�   -ZD  -8E  <W]  (8�  �   NY  D�-   Fe  >U   hY  H�"  $'$`  L�"  �"  �-  �-   QY  X?`  �-  �"  �"  �-   �Y  ]  �"  #  #  �-   yW  �uY  �"  +#  6#  �-  �"   X  ̄W  �"  N#  Y#  �-  �"   =�[  eoX  �"  	�"  y#  #  �-   =n\  l�\  �"  
�"  �#  �#  �-   =Z  t�X  �"  �"  �#  �#  �-  �"   =�W  ѲX  q  �"  �#   $  �-  �&  q   =P� ��^  �"  �"   $  +$  �-  �"   =�W  ��_  q  �"  K$  [$  �-  )  q   =� �:Z  N%  �"  {$  �$  �-   =09  �g^    �"  �$  �$  �-  z  �  �   ==H  �B_    �"  �$  �$  �-    �   >#`  �"  �$  %  �-  N%   	�"  !T  �%  ,�E  >     ?�  ?o  ?�  ?�  ?�  ?�  ?�	  @int ?(  ?#  ?�� ?�� ?�� :2*  7�%  A80    _� �2%  ?�  �  %  pW   +%  qW  !N%    "9%    #\%  BFd �%  .  <�%  `  DN%  �  W�%  �  _�%  �  eN%  t   mN%  a  uN%    ~N%  �  �N%  3  �N%  �  �N%  H  �N%  y  �N%    �N%  s  �N%  T   �N%  �  �N%  F  �N%  �  �N%  �  �N%    �N%  V  �N%  C�%  ?�  Ds  N�%  �  V�%  \	  2N%  o  7N%  �  <N%  �  CN%  �  N%  C�%  	\  �%  gX  �%  X\  &S'  X\  X,h(  $Z  .�%   \ /�%  � 1,'  Z  2�%  K]  3�%  �_  4�%  \W  5�%  �Z  6�%  -_  8�(   VY  9�(  $`  :�(  (�Y  ;�(  ,7_  <�(  0BY  = )  4b\  >�(  8\  ?�(  <7Y  @�(  @ Z  A1)  DSX  B1)  Hn4 D�%  L`  F�(  P*5 G�(  T E='  �(  �&  �%  �(   CS'  Ch(  E='  �(  �(  �%  �(   C�(  FC�(  EN%  �(  �(  2'  N%   C�(  E2'  �(  �(   C�(  EN%  �(  �(   C�(  E�(  )  )  )  �(   C)  	�%  C�(  G1)  �(   C&)  HpO qO !7)  IJ   Iz   ?�  Cz   CJ   I�  I�%  I)  C�   Iv"  Cv"  C�  I  ?  �  8�*  �{  �&   ]�  �&  \�   �&  �D  !�&  �3  "�&  U>  #�&  &�  $�&  �  %�&  �*  &�&   ڡ  '�%  $�U  (�%  %TL  )�%  &�I  *�%  'Q  +�%  (�C  ,�%  )�J  -�%  *1  .�&  ,o(  /�%  0�U  0�%  1PL  1�%  2�I  2�%  3Q  3�%  4�C  4�%  5�J  5�%  6 8)%  K�&  �*  N%  )   JGT  P�*  C�)  �    N%  	N%  CA  C�  C5  C.  I.  I�  I5  K2%  =+  L C�  I�  I�  �^  !!2'  MZ  !1l+  l+   CH'  8aY  !�N%  �+  l+   N\  !CN%  �+  l+   NxZ  !MN%  �+  l+   8`  !�N%  �+  l+   N�^  !rN%  �+  l+   N_X  !�N%  �+  l+  �+   CO+  N�_  !��&  ,  �&  N%  l+   8�\  !�l+  9,  )  )   N4Z  !��%  ^,  �(  �%  �%  l+   87`  !�l+  },  )  )  l+   N>]  !	N%  �,  l+  U%  N%   N�Z  !N%  �,  l+  �,   C�,  	O+  N�Y  ! U%  �,  l+   N�Y  !�N%  �,  l+   O\  !�N%  8�_  0�&  -  �&   M�]  !W"-  )   8D[  !TN%  7-  )   8�[  !aN%  Q-  )  )   M�\  !)c-  l+   PY@ !�y-  l+  �&   8�[  !�N%  �-  l+  �&  N%  �%   J�]  !il+  8D]  !w�&  �-  �&   N}W  !�N%  �-  N%  l+   C  Ca  I  Ia  	�-  Cf  C�"  Q�  .  .  Rh  .   	+  Q#  ,.  6.  Rh  .   C�  Q�  J.  ].  Rh  ].  R#  +   	6.  S�$  8r.  �.  Rh  �.  R#  +   	�-  T�  �.  U__c  �.   	P)  T�  �.  VhR  $�.  VmR  $�.   	i)  	i)  W�  T�  �.  U__c ,�.   	i)  C|  Q)  	/  /  Rh  /  U__c a�%   	�.  Q�"  2/  </  Rh  �.   Q#  J/  _/  Rh  �.  X__c Ǥ"   Q6#  m/  �/  Rh  �.  X__c ̤"   Q $  �/  �/  Rh  �.  X__c ��"  YZ�&  ��"    Q  �/  �/  Rh  .   Q  �/  �/  Rh  .   Q�  �/  �/  Rh  ].   QK  0  0  Rh  0  [Q  �z   	�-  Qf  00  :0  Rh  :0   	�-  I|  T�  d0  �R     X__f .�.   QZ  r0  �0  Rh  /  U__c 3�%   \d0  �T  ��   ��0  �0  ]r0  � ]{0  � \b.  X  `�   ��0  �0  ^r.  �Z  _<.  d�   8^J.  [  `v�  \b.  �W  ��$   �1  _1  ]r.  � ab.  ��   8U1  ^r.  0[  _<.  ��   8^J.  0[  b��  c���=   d#  ��   �v1  �1  eh  �.  � _$/  ��   o]2/  � f���,    dY#  ��    ��1  02  eh  �.  � g��   h__c g�"  O[  a$/  ��   g2  ]2/  � f���,   _</  ��   h]J/  � ^S/  O[  f���-     d�#  ��?   �G2  �2  eh  �.  � i__c t�"  �j�  k�&  v�"  b[  l�^  w%  _</  �   �^J/  u[  ^S/  �[  f��-     d[$  0�   ��2  �2  mh  �.  �[  c@��+   Q�$  �2  '3  Rh  �.  [Q  �z  [�J  ��  �  YZ�&  �  Z�_  �N%    \�2  g^  @�j   �B3  �3  ]�2  �]�2  �]�2  �]	3  �j�  n3  � o3  �[  a�/  \�   ��3  p0  ^0  �[   f��},  f���,    d+$  ��   ��3  �3  eh  �.  � i__s �)  �i__n �q  �f���=   d�#  ��M   �4  r4  eh  �.  � i__s ��&  �i__n �q  �j�  q�&  �q  Pa�.  ��   �g4  ^�.  �[   f��9,    \�/  �^   �I   ��4  5  ^�/  \  ^�/  .\  r�  �4  n�/  Ps_/  0��  �^m/  N\  ^v/  m\  cC�>    j   p�/  ^�/  �\  j   t�/  f[��+     u�$  p��   �5  �5  eh  �.  �v%  �  �v^F  ��  �w"0  }�  �a5  ]00  �� s�2  ��0  �^	3  �\  ^�2  �\  x�2  ^�2  �\  j0  t3  o3  �\  a�/  ��   ��5  ^0  ]  ^0  -]   f��},  f���,     y�   �   ��6  !T  �%  �E  >   �F  �  z%  �
�6  � z�^  �
�6  �{�/  �   �
y6  ]�/  �|.  �   �],.  �|.  �   -].  �   f�d    	C+  	&+  C%   Q�  �6  �6  Rh  �6  U__c ��%   	�6  }*    �s   ��7  !T  �%  �E  >   �F  �  z]\  �
�7  � z�^  �
�7  �~�6  +�H  �
�7  �6  
^�6  b]  ~E0  2�`  �R7  ^X0  �]  f���    ��.  6�x  �^/  �]  ^	/  �]  g`�.   ^/  �]  ^	/  ^  fi��     fN��    	I+  	,+  Q�"  �7  �7  Rh  �.  X__f L�-   \�7  \  ��Z   ��7  8  ]�7  � ]�7  �_�/  ��9   M^�/  ^  b��  d�"   �   �48  A8  eh  �.  �  �U  =N8   	�%  ��   >N8  �B  ?N8  ��  Ez8   	�%  �B   Fz8  �C  Gz8  �e  Hz8  �8  Iz8  ��  Jz8  �

  X�8   	�%  ��  Y�8  ��
  Z�8  l�   `�8  	�%  ��  f
9   	
&  ��  g
9  ��  h
9  ��  n69   	&  ��	  o69  ��  p69  �H  vb9   	 &  �`  wb9  �w  xb9  �   yb9  �~  �9   	+&  �   ��9  ��  ��9  �  ��9  ��   ��9  ��  ��9  ��	  ��9  ��  ��9   	6&  �  ��9  �  ��9  ��  ��9  ��  �4:   	A&  ��  �4:  ��  �4:  ��  �4:  �m  �m:   	L&  �	  �m:  �2	  �m:  ��  �m:  �9  �m:  �[  ��:   	W&  �J  ��:  ��  ��:  �7  ��:  ��  ��:   	b&  �I	  ��:  �$	  ��:  ��   �;   	m&  �N  �;  �p  �7;   	x&  ��  �7;  �:  �7;  ��  �7;  �d   �7;  ��  �};   	�&  �  �};  ��  �};  ��	  ѩ;   	�&  ��  ҩ;  �  ��;   	�&  ��  ��;  ��  ��;  ��  ��;  �+  �<   	�&  ��  �<  ��   �<  �  �-<   	�&  ��
  �-<  ��  �-<  �  �Y<   	�&  �   �Y<  �F  �Y<  ��  �<   	�&  ��  �<  ��  ��<  �D  O�<   	�&  ��  P�<  �1  Q�<  ��  W�<   	�&  �^  X�<  ��  3�<   	�&  ��  4�<  ��   8=   	 '  ��  9=  �l	  =:=  	'  �N  >:=  �^  ?:=  �L  @:=  �a  Ds=  	'  �B  Es=  ��	  Fs=  �  Gs=  �  Hs=  �y  Is=  ��   �=   	!'  ��  !�=  �  "�1  �=  �&   N�� !��%  >  �(  �%  �%  l+   �X  !�N%  N%  l+    �]   z   d  ib  �V  �-      �,  (  �  �  �  E   �  �  o  �	  �  qW  !s   int   "�   �  #  .  	<h   `  	Ds   �  	Wh   �  	_z   �  	es   t   	ms   a  	us     	~s   �  	�s   3  	�s   �  	�s   H  	�s   y  	�s     	�s   s  	�s   T   	�s   �  	�s   F  	�s   �  	�s   �  	�s     	�s   V  	�s   3   �  s  
N:   �  
V:   \	  2s   o  7s   �  <s   �  Cs   �  s   �  �  3   	pO qO !�  
std " 
)  @�  %  0�=  ��  �b  �3   Fe  �s   �3  �=  [  �*  �*   +  eq �<-  �*  }  �*  �*   lt ��1  �*  �  �*  �*   ��  eF  s   �  +  +  �   �K  �9  �  �  +   �(  
!  +  �  +  �  �*   1  �A  +     +  +  �   �5  �'  +  D  +  +  �   �3  �A  +  h  +  �  +   +  :  +  �  +   6  �C   �P  6  �  �*   �B  $6  �*  �  +  +   eof (�:  6  ?  ,N0  6  +    _� �,   5+  6E,  7_,  �?  �%   K  \�  *)   �e  _�  �4  c{,  �J  d�,  ��  qY  _  �,   ��  so  z  �,  �,   W  y�  �,  s       �J  p  �B  �     %  �   �B  �  �,  �  �,    �e  y%  [V  �  �  �G  !�   <  x  �4  {1  �J  |=  �J  �*  `S  ��*  ~J  �  �J  �  �%  ��  �K  ��   I  ��  :!  �p,   %H  �D  _    �3  2�   �G  7�   t3  B�,  !�'  ��O  �,  "V  ��N  �*  �  �  �,   "3  �o+  �*      �,   #�P  ��O    %  �,   #�M  ��P  8  >  �,   #�,  �-  Q  \  �,  �   "�+  ��R  �  s  y  �,   "3  �   �  �  �  �,  �,  �,   �/  !�B  �,  �  �  �  �,   #�O  �|6  �  �  �,  �,   $(  ��6  �    �,  �,   %�   �-  �      �,   &�1  o�*  �  3  �,  �,  �    %�A  $n%  �  \  b  �,   %�A  (�I  �  z  �  �,  �   %"A  ,�%  �,  �  �  �,   %�1  2E)  /  �  �  �,   %�/  6;&  /  �  �  �,   $�>  :�>  �  �  �,   %S  A:2  �    !  �,  �  �   $�#  K�(  5  J  �,  �  �  �   %9  S>$  �  b  r  �,  �  �   %-U  [�7  �*  �  �  �,  �   '�5  d�-  �  �  �  �   '	1  m�P  �  �  �  �   '�3  v\-  �  �  �  3    'nU  ��-  	  �  /  /   'nU  �nG  5	  �  ;  ;   'nU  ��   U	  �  �  �   'nU  �IP  u	  �  �  �   �J  �rR  s   �	  �  �   $�=  ��H  �	  �	  �,  �  �  �   $V  �)  �	  �	  �,   (�'  �D*  �,  )�0  ��	  �	  �,   *�0  �
  
  �,  �,   �0  �)
  4
  �,  �,   �0  �D
  Y
  �,  �,  �  �   �0  �i
  �
  �,  �,  �  �  �,   �0  ��
  �
  �,  �  �  �,   �0  ��
  �
  �,  �  �,   �0  ��
  �
  �,  �  3   �,   )�0  "�
  	  �,  s    +�  *,Q  �,  "  -  �,  �,   +�  2�G  �,  F  Q  �,  �   +�  =�%  �,  j  u  �,  3    +S� f�&  /  �  �  �,   +S� q�>  ;  �  �  �,   ,end y<  /  �  �  �,   ,end �6;  ;  �  �  �,   +I ��$  S  
    �,   +I ��7  G  )  /  �,   +��  �lC  S  H  N  �,   +��  �CM  G  g  m  �,   +r ��R  �  �  �  �,   +�K  �r5  �  �  �  �,   +�3  �j=  �  �  �  �,   -�� �  �  �  �,  �  3    -�� ��F      �,  �   +I  v  �  (  .  �,   -�E  �|U  C  N  �,  �   -�1  -�  c  i  �,   +�� 5�?  �*  �  �  �,   +�:  D�6  #  �  �  �,  �   +�:  UW    �  �  �,  �   ,at k
/  #  �  �  �,  �   ,at ��7        �,  �   +�F  ��/  �,  /  :  �,  �,   +�F  �k:  �,  S  ^  �,  �   +�F  ��H  �,  w  �  �,  3    +@  DA:  �,  �  �  �,  �,   +@  U�1  �,  �  �  �,  �,  �  �   +@  )�D  �,  �  �  �,  �  �   +@  ��*  �,    !  �,  �   +@  �6  �,  :  J  �,  �  3    -�G  -aN  _  j  �,  3    .�3  �b*  �,  �  �  �,  �,   +�3  ^ 2  �,  �  �  �,  �,  �  �   +�3  �=  �,  �  �  �,  �  �   +�3  z�T  �,  �    �,  �   +�3  � @  �,  !  1  �,  �  3    -� ��E  F  [  �,  /  �  3    +� �\+  �,  t  �  �,  �  �,   +� �u>  �,  �  �  �,  �  �,  �  �   +� g|=  �,  �  �  �,  �  �  �   +� "�@  �,  �    �,  �  �   +� 9k<  �,  '  <  �,  �  �  3    +� K�'  /  U  e  �,  /  3    +bL  d�R  �,  ~  �  �,  �  �   +bL  t�2  /  �  �  �,  /   +bL  �L&  /  �  �  �,  /  /   +�%  �9F  �,  �  	  �,  �  �  �,   +�%  �|<  �,  "  A  �,  �  �  �,  �  �   +�%  ��T  �,  Z  t  �,  �  �  �  �   +�%  ��A  �,  �  �  �,  �  �  �   +�%  b>  �,  �  �  �,  �  �  �  3    +�%  3%  �,  �    �,  /  /  �,   +�%  'V7  �,    6  �,  /  /  �  �   +�%  <�+  �,  O  d  �,  /  /  �   +�%  Q'S  �,  }  �  �,  /  /  �  3    +�%  vj.  �,  �  �  �,  /  /  �  �   +�%  ��9  �,  �  �  �,  /  /  �  �   +�%  �C  �,    0  �,  /  /  /  /   +�%  �>/  �,  I  c  �,  /  /  ;  ;   %�?  ��&  �,  {  �  �,  �  �  �  3    %�1  �O  �,  �  �  �,  �  �  �  �   ,)  �z-  �  �  �  3   �,   /+E  �3J  �    �  3   �,   +�5  ��)  �  '  <  �,  �  �  �   -n	 @D  Q  \  �,  �,   +W�  �6  �  u  {  �,   +�A  %�A  �  �  �  �,   +��  ,Z5    �  �  �,   +�(  �;  �  �  �  �,  �  �  �   +�(  I�%  �       �,  �,  �   +�(  X�5  �  )  9  �,  �  �   +�(  �^   �  R  b  �,  3   �   +�(  v�S  �  {  �  �,  �,  �   +�(  	K  �  �  �  �,  �  �  �   +�(  �o?  �  �  �  �,  �  �   +�(  J5  �  �    �,  3   �   +NW  ��Q  �  $  4  �,  �,  �   +NW  /�I  �  M  b  �,  �  �  �   +NW  ��,  �  {  �  �,  �  �   +NW  ��;  �  �  �  �,  3   �   +�S  ��I  �  �  �  �,  �,  �   +�S  >T?  �  �    �,  �  �  �   +�S  05  �  $  4  �,  �  �   +�S  $S:  �  M  ]  �,  3   �   +�>  2hL  �  v  �  �,  �,  �   +�>  SUB  �  �  �  �,  �  �  �   +�>  Q�2  �  �  �  �,  �  �   +�>  _�K  �  �    �,  3   �   +�4  qT  �    /  �,  �,  �   +�4  j�K  �  H  ]  �,  �  �  �   +�4  ��5  �  v  �  �,  �  �   +�4  N.  �  �  �  �,  3   �   +U+  �)  �  �  �  �,  �  �   +��  �!1  s   �  �  �,  �,   +��  ��T  s     *  �,  �  �  �,   +��  ��O  s   C  b  �,  �  �  �,  �  �   +��  �;.  s   {  �  �,  �   +��  ��B  s   �  �  �,  �  �  �   +��  ��,  s   �  �  �,  �  �  �  �   �  0!T  3   1�E    1�F     2�&  2�7  �  �o  >�   �| Cs   3Q  b<   #  3�F c<  3�R  d<  33  e<  3�  f<  3�K  g<  3�@  h<   4all i<  ?5�� ��  :!  �p,   NF  �&-  �E  ��  p0  �&-  �%  �2-  6S  �8-  6�R  �8-  63  �8-  6�$  �8-  6�K  �8-  6�@  �8-  6�@  �C-  $�4  �Z  S  Y  �,   $�=  y)  m  s  �,   7�� �  �  �,  Y-  �   7�� �  �  �,  �  �   7�� �  �  �,  �   7N  �  �  �,  s    7�� �    �,  Y-   $�  �U    #  �,  Y-   %�&  �.  �*  ;  A  �,   $�F  &�;  U  e  �,  _-  #   $�9  )�Q  y  �  �,  _-  N-   $WR  ,`2  �  �  �,  _-   -   $�S  /=  �  �  �,   -  ,-   8e  7,  �  �,  ,-  �    �$  �,   6OD  �,  6gP  �,  6�F  $�,  2< 9id ��  �U  ��   6�I  �p,  $�  �<?  b  m  -  -   :id �|  �  -  -   ;id ��  �  -   <4H  ��(  �  �   -    �o  u�  �  -   �o  ~�  �  -  -   *�o  ��    -  �   �o  �  *  -  -  �  #   �o  �:  O  -  -  -  #   5  �_  j  -  s    .�  ��*  -  �  �  -  -   .H�  ��N  �   �  �  -   .U  �9  �*  �  �  -  -   .2  �t*  �*  �  �  -  -   =jP  �D       -   >RD  �Q  -  ?�o  7-   8   -  �,   @�K  :�N  @�A  =�5  �K  @I  #  j   #   $�,  CH<  ~   �   -  -  -  #   (  #  �     � >�  AW  3B!  B�4  B�$  Bq-  Bc=  Bo'  B�5   B�%  � B�8  �BX)  �B�%  �B�  �BaO  �BY=  � BP  �� B�C  ��BwS  �B�O  � B�?  �B�5  �� A
$ g{!  B)W  B�   B�U  B�A  B�8  B�P   BEH  �� A�4  ��!  BO   B�7  B(  B�Q  BG  �� A��  ��!  B�R   B�-  B�1  BlO  �� Cb4 �#  D�  J{!  +l6 ��K  �'  �!  "  e1   +l6 �6N  �'  "  ("  �1  �'   +-H  ��`    A"  G"  e1   �P  ��   E�4  a"  G"  Fdec a"  Et-  a"  Fhex a"  Er'  a"  E< a"   Foct a"  @E� a"  �G[)  a"   G�%  "a"   G�  &a"   GdO  )a"   G\=  ,a"   G�P  /a"    G�C  3a"   @EzS  6a"  �E�O  9a"  JG�?  <a"  E�7  Nj#  �!  E(  Qj#  E�Q  Vj#  EO  Yj#   D�9  iB!  Fin w�#  �#  Fout z�#  D�N  ��!  Fcur ��#  �#   �a  $�$  rS  +a   Hm�  ,
$  �#  H��  -
$  H�4  .
$  H;�  /
$  H��  0
$  H� 1
$   H�� 2
$  @Ib  3
$  I�e  4
$   I�  5
$   Hމ  6
$   �!  C�Y  �%  5�_ ��$  �M  ��*   *�_ .�$  �$  j-  p-  �*   <�  ��e  �*  �$  v-    b  J�&  �$  .�d  %�c  p-  %  .%  �3  �3  �'  .%   �b  >3   Fe  ?6  :%  {'  E�%  .%  .Ic  pb  p-  t%  �%  �3  �'  :%   0!T  3   1�E    <Ic  o�d  p-  �%  �3  �'    C�M  �&  +�* �e  �-  �%  �%  �-   �b  �3   +�* �_e  �-  &  
&  �-   -\b  (a  &  *&  |-  �'   -cb  �Pc  ?&  J&  |-  s    +�a  R(b  i&  c&  i&  |-   Fe  �6  +�c  <�c  i&  �&  �&  |-   +!a  *�a  i&  �&  �&  |-   0!T  3   1�E     C�+   '  Jis 1�c  �*  �&  �&  �1  �#  3    KOe  ��c  �  
'  �1  �#  �  �    C�E  �'  +3F  ;�S  |-  B'  H'  �-   .9U  ؍0  �!  `'  f'  �-   .�M  ��B  �!  ~'  �'  �-   LeU  ��4  �'  �'  �2  �!   LbU  �IQ  �'  �'  �2  �!   0!T  3   1�E    M�1  )�%  �'  �2  �!     '  �%  �>  b  N�*  �{!  (  {!  {!   N	W  �1  9(  1  {!   {!  N*  �{!  X(  {!  {!   �&  �  N�b  2  �(  O_Tp %   �2  �2   /c  �da  p-  �(  p-  �   �`  �b  p-  �(  p-  �,   �'  t\  e�Z  p-  �(  p-  �,  3    P}`  ��d  �]  0�R  �&  -    Q$   ��*  �  $,�  -  K  :�*  �e  =�  � ?�  "  @�  �4  A{,  �J  B�,  �A  O�)  �)  �,   �A  Q�)  �)  �,  �,   �A  V�)  �)  �,  s    .�
 Y51  B)  �)  �)  �,  Z)   .�
 ]�R  N)  �)  *  �,  f)   .� c?  B)  *  ,*  �,  6)  �   L_ m.   @*  P*  �,  B)  6)   .�3  q89  6)  h*  n*  �,   L.E  ��3  �*  �*  �,  B)  �,   L�(  ��(  �*  �*  �,  B)   O_Tp 3    *)  2ZD  28E   �� �� �� Q2*  7�*  R8   S+  S[  �  [  +  S�  �  8 E,  �{   �   ]�   �  \�    �  �D   !�  �3   "�  U>   #�  &�   $�  �   %�  �*   &�   ڡ   '3   $�U   (3   %TL   )3   &�I   *3   'Q   +3   (�C   ,3   )�J   -3   *1   .�  ,o(   /3   0�U   03   1PL   13   2�I   23   3Q   33   4�C   43   5�J   53   6 N)%   K�  _,  s   �   TGT   Pj,  +  �  ! s   S3   S�  *)  S�*  �*    S�    �*  �    �  �  S�  S  S�  U,   �,  V �  �  �,  �,  �    S�   �   (  S�   �   ,-  �   �  U -  C-  V UN-  N-  V T-   -  S�   �   %   �$  S�$  �$  �%  �'  W)'  �-  �-  Xh  �-   �-  �%  �'  W�%  �-  �-  Xh  �-   �-  W�%  �-  �-  Xh  �-   W
&  �-  
.  Xh  
.  Y__n �'   |-  W�  .  '.  Xh  '.   �,  W*&  :.  P.  Xh  
.  Y__n �s    WH'  ^.  h.  Xh  �-   Wf'  v.  �.  Xh  �-   W�  �.  �.  Xh  �.   �,  WD  �.  �.  Xh  '.   W�  �.  �.  Xh  '.   Wm  �.  �.  Xh  '.   W%  �.  �.  Xh  �.   �,  WJ  /  @/  Xh  '.  Z%  S�  ZQ  S�  [\�c  U�,    W�  N/  p/  Xh  '.  Z%  A�  Y__s A�   ]A  �/  ^hR  �/  ^mR  �/   �*  �*  ]�  �/  [___p ��    W\  �/  �/  Xh  �.   W>  �/  �/  Xh  �.  `__n ��   W  �/  0  Xh  '.   ]�  50  Y__s 
+  Y__n 
�  Y__a 
50   �*  ]h  Q0  Y__c Q0   +  ]�  m0  Y__c  m0   �*  WJ&  �0  �0  Xh  
.  [\�&  Ti&    Wu&  �0  �0  Xh  
.  [\�&  >i&    ]�  �0  ZhR  $�0  ZmR  $�0   +  +  a�  ](  1  `__a �{!  `__b �{!   S9(  S{!  ](  ?1  `__a �?1  `__b �{!   1  ]>(  e1  `__a �{!  `__b �{!   �$  W�!  y1  �1  Xh  �1   e1  �!  W"  �1  �1  Xh  �1  Z�R  ��'  [\'U  ��'    �1  X(  W�&  �1  62  Xh  62  `__m 2�#  `__c 23   [b�&  8�*  b�`  9](  b�b  :�  [ba  =
$  [b�c  @�*      �1  W�&  I2  t2  Xh  62  `__m ��#  ^�a  ��  ^�a  ��   W�$  �2  �2  Xh  �2   v-  Se-  ]b(  �2  O_Tp %   `__a ��2  `__b ��2   �2  �2  ]   �2  Z�e  +  Z�e  +  Y__n �    '  W�'  3  #3  Xh  #3  ^�%  ��!   �2  W�'  63  K3  Xh  #3  ^�%  ��!   W("  Y3  c3  Xh  �1   W^  q3  �3  Xh  �3  Y__c �3    �,  W�&  �3  �3  Xh  
.  [\�&  ,i&    �$  .%  c%  �  ��3  �9  dh  �9  � e__s &�3  4^  f__n &�'  �g�e  &.%  �h  �9  i�*  )�!  _  j�$  *�$  �_h@  �7  i�a  /F%  ]_  i�^  0F%  �_  i(  1�9  �_  k__c 2:%  `  lV0  ?�   /�4  m`0  *`   nr0  S�h  2 5  m�0  �_  oS�   �4  p�0  qV0  _�   Vm`0  �`    r_�!   m�0  �`  r_�!   p�0     h�  L7  i�a  8�'  �`  h�  '6  ___p >�9  n0  b��  @d5  m(0  a  m0  Ma  m0  ka  s���\   n�2  ���  C�5  m�2  �`  m�2  ~a  m�2  �a  s�� ]   n�-  ��   E�5  m�-  �a  m�-  �a   tr0  ��0   Gm�0  b  hX   6  p�0  qV0  	�   Vm`0  :b    r �    m�0  Yb  r �    p�0      n:0  ��x   KD6  mD0  xb   t�3  ���   Mm�3  �b  u�   v�3  c  w�0  ���   .�6  m�0  �b  o��
   �6  v�0  Jc  q,.  ��   Bx:.  mC.  hc    r@�   m�0  |c  r@�   p�0     yr0  ��   /m�0  �c  o�
   &7  p�0  qV0  �   Vm`0  �c    r��   m�0  �c  r��   p�0        l1  ��   Yj7  x31  x(1   n�0  ���   V�7  m�0  �c  h !  �7  p�0  y,.  ��!  Bx:.  mC.  $d    r��   m�0  8d  r��   p�0     z1  ��   Rx31  x(1    n(3  �0!  ai8  m?3  Wd  m63  wd  l1  $�   �_8  m31  Wd  m(1  �d  z�0  $�   �m1  Wd  m�0  �d    s�>]   hP!  
9  {�9  n(3  ��h!  ]�8  m?3  �d  m63  �d  l1  ��   ��8  m31  �d  m(1  	e  z�0  ��   �m1  �d  m�0  +e    s��>]   s��D]  s��X]  s��>]   l1  d�   h09  m31  ?e  m(1  Se   n 3  i��!  j�9  m3  ke  m3  ~e  l�0  q�   �{9  m1  ke  m�0  �e   s{��'   |2�s�D]  s7�X]  s�X]   s��^]  s�^]   �3  K%  W%  Q  " �9  2�  �9  S�9  c\%   ��  ��9  ?  dh  �9  � f__n q�'  �g�e  q:%  �h�!  ?  j�$  w�$  �_h�!  �>  i�*  z�!  �e  h�!  l=  ia  }W%  �e  i�^  ~F%  7f  i(  �9  ff  k__c �:%  �f  iAc  ��*  g  l:0  j�   }�:  mD0  Ag   nr0  � "  �1;  m�0  ff  o�   ;  p�0  qV0  ��   Vm`0  yg    rf�   m�0  �g  rf�   p�0     h"  �<  i�a  ��'  �g  h@"  �;  ___p ��9  n0  ��`"  ��;  m(0  �g  m0  �g  m0  �g  s���\   nr0  ���"  ��;  m�0  �g  u�"  p�0  qV0  �   Vm`0  h     t�-  ���"  �m�-  h  m�-  �g    t�3  ���"  �m�3  ,h  u�"  v�3  Xh  w�0  ���"  .�<  m�0  ,h  h#  o<  v�0  �h  q,.  ��	   Bx:.  mC.  �h    r�   m�0  �h  r�   p�0     qr0  ��0   /m�0  �h  o��   �<  p�0  qV0  ��   Vm`0  �h    r��   m�0  �h  r��   p�0        t�0  �(#  �m�0  i  o�   H=  p�0  q,.  �   Bx:.  mC.  >i    rz�!   m�0  Ri  rz�!   p�0      n 3  R�@#  ��=  m3  fi  m3  zi  l�0  Q�   ��=  m1  fi  m�0  �i   s^��'   h`#  b>  {?  n(3  ��x#  �F>  m?3  �i  m63  �i  l1  ��   �<>  m31  �i  m(1  �i  z�0  ��   �m1  �i  m�0  j    s��>]   s��D]  s��X]  s�>]   n(3  ���#  ��>  m?3  j  m63  5j  l1  ��   ��>  m31  j  m(1  Sj  z�0  ��   �m1  j  m�0  uj    s�>]   s��D]  s��X]  s�X]   |L�s���%   s��^]  s�^]   �9  }�(   ��  �:F  ge  �:F  � e__s Ņ  �j  h�#  'F  De  �:%  {'  �K%  b  ��$  i�d  ��'  k  i�*  ��!  �k  j�$  Й$  �[h�#  �D  i	e  ��'  �k  i�b  ��?  'l  �?  S�?  k?  i�^  ��?  ^l  U?  i(  ��?  �l  `?  k__c �U?  �l  nK3  J� $  �/@  xY3  |q� nr0  �� $  ޗ@  m�0  �l  h@$  t@  p�0  qV0  ��   Vm`0  &m    r|�"   m�0  9m  r|�"   p�0     hX$  �C  i�a  ��'  Mm  n;2  '��$  �A  mh2  km  m]2  �m  mR2  �m  mI2  4n  u�$  xh2  m]2  ln  xR2  xI2  t�1  ���$  �m�1  �n  m�1  �n  m�1  o  u�$  m�1  o  m�1  �n  m�1  �n  u�$  v�1  0o  p2  v2  ho  u%  v2  p  u8%  v'2  p  s��r]  s2��]  s���]  s���]  s��]         l�2  v�   ��A  m�2  Mm  m�2  �p  m�2  �p  s�� ]   n�-  ��h%  �B  m�-  �p  m�-  q   nr0  ���%  �B  m�0  �p  h�%  \B  p�0  qV0  ��   Vm`0  -q    r0�   m�0  Lq  r0�   p�0     t�3  )��%  �m�3  `q  u�%  v�3  �q  w�0  )� &  .C  m�0  `q  o)�   �B  v�0  �q  q,.  1�   Bx:.  mC.  �q    rD�   m�0  �q  rD�   p�0     yr0  7�&  /m�0  #r  o7�   aC  p�0  qV0  ?�   Vm`0  Cr    re�   m�0  Vr  re�   p�0        n�1  ��0&  �3D  m�1  jr  m�1  �r  m�1  s  uX&  x�1  x�1  x�1  uX&  v�1  ms  p2  v2  �s  up&  v2  t  u�&  v'2  �t  s��r]  s���]  sl��]  s���]  s���]       l:0  ��   �PD  mD0  u   w�1  ���&  �D  m�1  Xu  m�1  �u  u�&  v�1  �u    sy��(  |��|�� w(3  ���&  E  m?3  �u  m63  v  l1  ��   �E  m31  �u  m(1  ,v  z�0  ��   �m1  �u  m�0  Nv    s�>]   o��=   �E  {?F  w(3  ���&  �E  m?3  bv  m63  vv  l1  ��   ��E  m31  bv  m(1  �v  z�0  ��   �m1  bv  m�0  �v    s��>]   s��D]  s��X]  s��>]   ~ 3   �   F  x3  m3  �v  l�0  #�   ��E  x1  m�0  �v   s-��'   |7�s��D]  s	�X]  s�X]   s��^]  s�^]   p-  �9  We  RF  tF  Xh  �3  Z%  d�  Y__n d�   WJ  �F  �F  Xh  �3  Y__c -3   [\R'  /�    }�(   �X  ��O  e  �O  � �^  �O  �h'  �O  �De  :%  �{'  K%  �b  �$  ��e  �  ��d   G  �v  ��*  !�!  Ew  ��$  "�$  �[h0'  �M  �__w (�(  �__n )mG  �w  G  ��b  +�G  �w  �G  S�G  �F  ��^  ,�G  �w  �F  �(  -�G  �w  �F  �__c .�F  Lx  wDF  {�h'  'YH  �gF  �[F   mRF  �x  w/  {��'  gOH  �%/  �/   m/  �x  u�'  �2/   y�.  {��'  Um�.  �x     s���	   wK3  ���'  +xH  xY3  |�� wr0  ���'  .�H  m�0  �w  h�'  �H  p�0  qV0  ��   Vm`0  �x    u�'  m�0  �x  u�'  p�0     h�'  �L  ��a  5�'  �x  w�3  ��8(  G�I  m�3  y  u8(  v�3  Ey  w�0  ��`(  .�I  m�0  y  h�(  mI  v�0  ty  y,.  ���(  Bx:.  mC.  �y    rL�   m�0  �y  rL�   p�0     yr0  ���(  /m�0  �y  h�(  �I  p�0  qV0  ��   Vm`0  �y    r&�   m�0  �y  r&�   p�0       w;2  Q��(  <K  mh2   z  m]2  4z  mR2  �z  mI2  �z  u)  xh2  m]2  {  xR2  xI2  t�1  0�0)  �m�1  *{  m�1  j{  m�1  �{  u0)  m�1  �{  m�1  *{  m�1  j{  u0)  v�1  �{  p2  v2  �{  uX)  v2  �|  u�)  v'2  }  s|�r]  sR��]  s���]  s��]  s<��]         w�-  ���)  ?)K  m�-  S}  m�-  f}   wr0  ���)  ARK  m�0  y}  u�)  p�0    wc3  ���)  E�L  mz3  �}  mq3  �}  ytF  ���)  �m�F  �}  m�F  �}  u�)  v�F  �}  ~�.  ��   /�K  m�.  �}  q�.  ��   �m�.  �}  q�.  ��   -m�.  �}     ~p/  ��   2!L  m�/  �}  mz/  %~   ~�.  ��   3YL  m�.  =~  q�.  ��   -m�.  =~    w�/  ��*  3�L  m�/  i~  m�/  �~  r��   m�/  �~  m�/  �~  l�.  ��   ճL  x�.   zp/  ��	   �x�/  mz/  �~     s��.     s���   w�1   � *  3�M  m�1  �~  m�1  _  m�1  �  uH*  x�1  x�1  x�1  uH*  v�1  �  p2  v2  �  u`*  v2  i�  u�*  v'2  )�  s��r]  s���]  s���]  s���]  s���]       ~:0  �   3�M  mD0  s�   w�1  ���*  M�M  m�1  ��  m�1  �  u�*  v�1  B�    s���(  |��|�� h�*  �N  {�O  w(3  ���*  Q�N  m?3  ��  m63  ��  l1  ��   �zN  m31  ��  m(1  ��  z�0  ��   �m1  ��  m�0  ��    s��>]   s��D]  s�X]  s-�>]   w(3  <�+  YO  �?3  m63  �  l1  D�   �O  �31  m(1  �  z�0  D�   ��1  m�0  4�    sh�>]   ~ 3  V�   _`O  x3  m3  H�  l�0  Y�   �VO  x1  m�0  [�   sc��'   |7�s6�D]  sS�X]  so�X]   s(�^]  sx�^]   p-  �,  �9  }�(  ��  �WW  e  eWW  � �^  e\W  ��e  f3   �h(+  DW  �De  i:%  ��b  j.%  �{'  lK%  ��e  n�  ��d  pP  o�  �__n qBP  ���?P  ��*  r�!  �  ��$  s�$  �_hH+  �U  ��a  y�P  H�  �O  ��^  z�P  ��  �(  {�P  ��  P  �__c |�O  ��  hx+  5T  \�a  ��'  w�3  ���+  ��Q  m�3  -�  u�+  v�3  V�  wr0  ���+  /iQ  m�0  ��  h�+  FQ  p�0  qV0  ��   Vm`0  ��    r@�   m�0  ��  r@�   p�0     y�0  #�,  .m�0  -�  o#�
   �Q  v�0  ��  q,.  '�   Bx:.  mC.  ܅    r��   m�0  ��  r��   p�0       h ,  �R  �__p ��Q  �Q  �O  w0  �@,  �7R  m(0  �  m0  &�  m0  E�  sW��\   w�-  q�h,  �ZR  m�-  d�  x�-   wr0  {��,  ��R  m�0  w�  u�,  p�0    sq��   ~:0  ��   ��R  mD0  ��   yc3  ���,  �mz3    mq3  ׆  ytF  ���,  �m�F    m�F  ׆  u�,  v�F  �  ~�.  ��   /OS  m�.  ׆  q�.  ��   �m�.  ׆  q�.  ��   -m�.  ׆     ~p/  �   2vS  m�/  "�  mz/  J�   ~�.  
�   3�S  m�.  b�  q�.  
�   -m�.  b�    w�/  ��,  3(T  m�/  ��  m�/  ��  r��   m�/  ܇  m�/  ��  l�.  ��   �T  x�.   zp/  ��	   �x�/  mz/  �     s��.      wDF  ���,  x�T  �gF  �[F   mRF  �  w/  ���,  g�T  �%/  �/   m/  �  u�,  �2/   y�.  ���,  Um�.  �     s���	   ~V0  ��   y�T  m`0  V�   wr0  �-  |HU  m�0  ��  o�   %U  p�0  qV0  
�   Vm`0  ҈    r��   m�0  �  r��   p�0     y�0  �� -  �m�0  �  o��   �U  p�0  q,.  ��   Bx:.  mC.  !�    r��   m�0  5�  r��   p�0      o�=   ]V  {aW  w(3  �8-  �AV  m?3  H�  m63  h�  l1  �   �7V  m31  H�  m(1  ��  z�0  �   �m1  H�  m�0  ��    s,�>]   s�D]  s5�X]  sC�>]   w(3  R�P-  ��V  m?3  ��  m63  ܉  l1  Z�   ��V  m31  ��  m(1  ��  z�0  Z�   �m1  ��  m�0  �    s��>]   w 3  ��p-  �#W  x3  m3  0�  l�0  ��   �W  x1  m�0  C�   s���'   |��sL�D]  si�X]  s��X]   s>�^]  s��^]   p-  �,  �9  �U  	=sW   �   ��   	>sW  �B  	?sW  ��  	E�W   �   �B   	F�W  �C  	G�W  �e  	H�W  �8  	I�W  ��  	J�W  �

  	X�W   �   ��  	Y�W  ��
  	Z�W  ��   	`X  �   ��  	f0X   �   ��  	g0X  ��  	h0X  ��  	n\X   �   ��	  	o\X  ��  	p\X  �H  	v�X   �   �`  	w�X  �w  	x�X  �   	y�X  �~  	�X   �   �   	��X  ��  	��X  �  	��X  ��   	��X  ��  	��X  ��	  	��X  ��  	�!Y   �   �  	�!Y  �  	�!Y  ��  	�!Y  ��  	�ZY   �   ��  	�ZY  ��  	�ZY  ��  	�ZY  �m  	��Y     �	  	��Y  �2	  	��Y  ��  	��Y  �9  	��Y  �[  	��Y     �J  	��Y  ��  	��Y  �7  	��Y  ��  	�Z     �I	  	�Z  �$	  	�Z  ��   	�>Z   "  �N  	�>Z  �p  	�]Z   -  ��  	�]Z  �:  	�]Z  ��  	�]Z  �d   	�]Z  ��  	ɣZ   8  �  	ʣZ  ��  	ˣZ  ��	  	��Z   C  ��  	��Z  �  	��Z   N  ��  	��Z  ��  	��Z  ��  	��Z  �+  	�'[   Y  ��  	�'[  ��   	�'[  �  	�S[   d  ��
  	�S[  ��  	�S[  �  	�[   o  �   	�[  �F  	�[  ��  	�[   z  ��  	��[  ��  	��[  �D  
O�[   �  ��  
P�[  �1  
Q�[  ��  
W\   �  �^  
X\  ��  3"\   �  ��  4"\  ��   8A\   �  ��  9A\  �l	  =`\  �  �N  >`\  �^  ?`\  �L  @`\  �a  D�\  �  �B  E�\  ��	  F�\  �  G�\  �  H�\  �y  I�\  ��   �\   �  ��  !�\  ��`  �`  �   ]  �  s   ,    ��d  �  >]  �  �  �   ��  ��  �  X]  �   ��  �>  Y  r]  �   N�e  #rs   �]  s    Nb  #^s   �]  s    N�e  #Js   �]  s    NWe  #|s   �]  s    N�d  #�s   �]  s    SX(   ]g  �(   �  Bn  �V  �      �:  (  _� �7   �  �  8k  �{  k   ]�  k  \�   k  �D  !k  �3  "k  U>  #k  &�  $k  �  %k  �*  &k   ڡ  'q  $�U  (q  %TL  )q  &�I  *q  'Q  +q  (�C  ,q  )�J  -q  *1  .k  ,o(  /q  0�U  0q  1PL  1q  2�I  2q  3Q  3q  4�C  4q  5�J  5q  6 q  �  std 2 �j  5>   6�j  7�j  @�l  	++ S	��  Y	%+  \�$ _�  
�    ��  c�  
�    �  g�  
�    %  *0a1  v!  �#  �  _Tp �.  �?  �    �=  ��  �b  �q  Fe  �j  �3  �=  ]  �t  �t   -  eq �<-  �t    �t  �t   lt ��1  �t  �  �t  �t   ��  eF  �j  �  �t  �t  �   �K  �9  �  �  �t   �(  
!  �t  �  �t  �  �t   1  �A  �t  "  �t  �t  �   �5  �'  �t  F  �t  �t  �   �3  �A  �t  j  �t  �  -   +  :  -  �  �t   8  �C   �P  8  �  �t   �B  $6  �t  �  �t  �t   eof (�:  8  ?  ,N0  8  �t    _� �7   �?  �%   K  \  �l   �e  _�  �4  c�t  �J  d�t  ��  qF  L  �t   ��  s\  g  �t  �t   W  ys  �t  �j    �  �J  	p�  �B  	�  
�   %  	k   �B  	�  �  u  k  �t   �B  �  u  �j    �e  	y   [V  	�  �  �G  	!�   <  	x�  �4  	{  �J  	|*  �J  	n  `S  	��p  ~J  	��  �J  	��  �%  	��  �K  	��   I  	��  :!  	��t   %H  	�I  
d   !�3  2�  !�G  7�j  !t3  B0u  "�'  	��O  u  #V  	��N  �t  �  �  ;u   #3  	�o+  �t      ;u   $�P  	��O  $  *  u   $�M  	��P  =  C  u   $�,  	�-  V  a  u  �   #�+  	��R  k  x  ~  u   #3  	�   k  �  �  u  �t  �t   �/  !�B  u  �  �  �  �t   $�O  	�|6  �  �  u  �t   %(  ��6  �    u  �t   &�   	�-  k    $  u   '�1  o�*  k  8  u  �t  �    &�A  	$n%  k  a  g  u   &�A  	(�I  k    �  u  k   &"A  	,�%  u  �  �  u   &�1  	2E)  4  �  �  u   &�/  	6;&  4  �  �  u   %�>  	:�>  �  �  u   &S  	A:2  �    &  u  �  �j   %�#  	K�(  :  O  u  �  �  �j   &9  	S>$  �  g  w  u  �  �   &-U  	[�7  �t  �  �  u  �j   (�5  	d�-  �  k  �j  �   (	1  	m�P  �  k  �j  �   (�3  	v\-  �  k  �  q   (nU  	��-  	  k  4  4   (nU  	�nG  :	  k  @  @   (nU  	��   Z	  k  k  k   (nU  	�IP  z	  k  �j  �j   �J  	�rR  �j  �	  �  �   %�=  ��H  �	  �	  u  �  �  �   %V  �)  �	  �	  u   )�'  	�D*  u  *�0  	��	  
  u   +�0  �
  
  u  �t   �0  �.
  9
  u  $u   �0  �I
  ^
  u  $u  �  �   �0  �n
  �
  u  $u  �  �  �t   �0  ��
  �
  u  �j  �  �t   �0  ��
  �
  u  �j  �t   �0  ��
  �
  u  �  q  �t   *�0  	"    u  �j   ,�  	*,Q  *u  '  2  u  $u   ,�  	2�G  *u  K  V  u  �j   ,�  	=�%  *u  o  z  u  q   ,S� 	f�&  4  �  �  u   ,S� 	q�>  @  �  �  u   -end 	y<  4  �  �  u   -end 	�6;  @  �  �  u   ,I 	��$  X      u   ,I 	��7  L  .  4  u   ,��  	�lC  X  M  S  u   ,��  	�CM  L  l  r  u   ,r 	��R  �  �  �  u   ,�K  	�r5  �  �  �  u   ,�3  	�j=  �  �  �  u   .�� �  �  �  u  �  q   .�� 	��F  	    u  �   ,I  	v  �  -  3  u   .�E  �|U  H  S  u  �   .�1  	-�  h  n  u   ,�� 	5�?  �t  �  �  u   ,�:  	D�6  (  �  �  u  �   ,�:  	UW    �  �  u  �   -at 	k
/  (  �  �  u  �   -at 	��7        u  �   ,�F  	��/  *u  4  ?  u  $u   ,�F  	�k:  *u  X  c  u  �j   ,�F  	��H  *u  |  �  u  q   ,@  DA:  *u  �  �  u  $u   ,@  U�1  *u  �  �  u  $u  �  �   ,@  )�D  *u  �    u  �j  �   ,@  	��*  *u    &  u  �j   ,@  �6  *u  ?  O  u  �  q   .�G  	-aN  d  o  u  q   /�3  �b*  *u  �  �  u  $u   ,�3  	^ 2  *u  �  �  u  $u  �  �   ,�3  �=  *u  �  �  u  �j  �   ,�3  	z�T  *u      u  �j   ,�3  	� @  *u  &  6  u  �  q   .� 	��E  K  `  u  4  �  q   ,� 	�\+  *u  y  �  u  �  $u   ,� 	�u>  *u  �  �  u  �  $u  �  �   ,� g|=  *u  �  �  u  �  �j  �   ,� 	"�@  *u      u  �  �j   ,� 	9k<  *u  ,  A  u  �  �  q   ,� 	K�'  4  Z  j  u  4  q   ,bL  	d�R  *u  �  �  u  �  �   ,bL  	t�2  4  �  �  u  4   ,bL  �L&  4  �  �  u  4  4   ,�%  	�9F  *u  �    u  �  �  $u   ,�%  	�|<  *u  '  F  u  �  �  $u  �  �   ,�%  ��T  *u  _  y  u  �  �  �j  �   ,�%  	��A  *u  �  �  u  �  �  �j   ,�%  	b>  *u  �  �  u  �  �  �  q   ,�%  	3%  *u  �    u  4  4  $u   ,�%  	'V7  *u  !  ;  u  4  4  �j  �   ,�%  	<�+  *u  T  i  u  4  4  �j   ,�%  	Q'S  *u  �  �  u  4  4  �  q   ,�%  	vj.  *u  �  �  u  4  4  k  k   ,�%  	��9  *u  �    u  4  4  �j  �j   ,�%  	�C  *u    5  u  4  4  4  4   ,�%  	�>/  *u  N  h  u  4  4  @  @   &�?  ��&  *u  �  �  u  �  �  �  q   &�1  �O  *u  �  �  u  �  �  �j  �   ,)  	�z-  k  �  �  q  �t   0+E  �3J  k    �  q  �t   ,�5  ��)  �  ,  A  u  k  �  �   .n	 @D  V  a  u  *u   ,W�  	�6  �j  z  �  u   ,�A  	%�A  �j  �  �  u   ,��  	,Z5    �  �  u   ,�(  �;  �  �  �  u  �j  �  �   ,�(  	I�%  �      u  $u  �   ,�(  	X�5  �  .  >  u  �j  �   ,�(  �^   �  W  g  u  q  �   ,�(  	v�S  �  �  �  u  $u  �   ,�(  	K  �  �  �  u  �j  �  �   ,�(  	�o?  �  �  �  u  �j  �   ,�(  J5  �       u  q  �   ,NW  	��Q  �  )  9  u  $u  �   ,NW  /�I  �  R  g  u  �j  �  �   ,NW  	��,  �  �  �  u  �j  �   ,NW  	��;  �  �  �  u  q  �   ,�S  	��I  �  �  �  u  $u  �   ,�S  >T?  �  �    u  �j  �  �   ,�S  	05  �  )  9  u  �j  �   ,�S  	$S:  �  R  b  u  q  �   ,�>  	2hL  �  {  �  u  $u  �   ,�>  SUB  �  �  �  u  �j  �  �   ,�>  	Q�2  �  �  �  u  �j  �   ,�>  _�K  �  �    u  q  �   ,�4  	qT  �  $  4  u  $u  �   ,�4  j�K  �  M  b  u  �j  �  �   ,�4  	��5  �  {  �  u  �j  �   ,�4  N.  �  �  �  u  q  �   ,U+  	�)  �  �  �  u  �  �   ,��  	�!1  �j  �    u  $u   ,��  ��T  �j    /  u  �  �  $u   ,��  ��O  �j  H  g  u  �  �  $u  �  �   ,��  �;.  �j  �  �  u  �j   ,��  ��B  �j  �  �  u  �  �  �j   ,��  ��,  �j  �  �  u  �  �  �j  �   �  0<�  { �  k  "  ß  �j  �j  �j  �t  �   ��  	���  k  T  �  �j  �j  �j  �t  �   <�  	�Ģ  k  �  �  �j  �j  �j  �t   �  ��  �  f�  �j  u  �j  �j  �t   !T  q  1�E  !  1�F  �   2�&  2�7  �  �o  >�!  �| C�j  3Q  b�   �  3�F c�  3�R  d�  33  e�  3�  f�  3�K  g�  3�@  h�   4all i�  ?5�� ��  :!  ��t   NF  �{u  �E  ��  p0  �{u  �%  ��u  6S  ��u  6�R  ��u  63  ��u  6�$  ��u  6�K  ��u  6�@  ��u  6�@  ��u  %�4  �Z      Au   %�=  y)  0  6  Au   �� F  V  Au  �u  �   �� f  v  Au  �j  �   �� �  �  Au  �   N  �  �  Au  �j   �� �  �  Au  �u   %�  �U  �  �  Au  �u   &�&  �.  �t  �    Au   %�F  &�;    (  Au  �u  �   %�9  )�Q  <  L  Au  �u  �u   %WR  ,`2  `  p  Au  �u  uu   %�S  /=  �  �  Au  uu  �u   7e  7,  �  Au  �u  �    �$  Au   6OD  Au  6gP  Au  6�F  $Gu  8< }  9< r     ��  �   :�h  �ܧ  "  Ae  ;��  ���  �j  :��  z�r  T  Ae �j  �-   ;�m  �~�  �-  <��  ~�  �-  Ae   =id �   �U  ��   6�I  ��t  %�  �<?  �  �  iu  ou   >id ��  �  iu  ou   ?id ��  �  iu   @4H  ��(  �     uu    �o  u   $   Wu   �o  ~4   ?   Wu  ]u   +�o  �O   Z   Wu  �j   �o  �j      Wu  ]u  �j  �   �o  ��   �   Wu  ]u  ]u  �   5  ��   �   Wu  �j   /�  ��*  ]u  �   �   Wu  ]u   /H�  ��N  �!  �    !  cu   /U  �9  �t  !  #!  cu  ]u   /2  �t*  �t  ;!  F!  cu  ]u   AjP  �D  �  a!  ]u   ;RD  �Q  ]u  B�o  7�!  �!  Wu  Au   C�K  :�N  C�A  =�5  �K  @I  �  �!  �   %�,  CH<  �!  �!  Wu  ]u  ]u  �   }  �  _   �  � >�  �a  $�"  rS  +k  Dm�  ,+"  "  D��  -+"  D�4  .+"  D;�  /+"  D��  0+"  D� 1+"   D�� 2+"  @Eb  3+"  E�e  4+"   E�  5+"   Dމ  6+"   FW  3;#  G�4  G�$  Gq-  Gc=  Go'  G�5   G�%  � G�8  �GX)  �G�%  �G�  �GaO  �GY=  � GP  �� G�C  ��GwS  �G�O  � G�?  �G�5  �� F
$ gt#  G)W  G�   G�U  G�A  G�8  G�P   GEH  �� F�4  ��#  GO   G�7  G(  G�Q  GG  �� 8b4 &  H�  Jt#  ,n4 '�T  �#  �#  �#  �   �P  ��"  ,n4 2�t  �#  �#  $  7�  �#   ,�/ m��  /M  $  %$  �   ,l6 ��K  /M  >$  D$  �   ,l6 �6N  /M  ]$  h$  7�  /M   ,*H  ��7  ]u  �$  �$  �   ,-H  ��`  �  �$  �$  �   �#  I�4  �$  Jdec �$  It-  �$  Jhex �$  Ir'  �$  I< �$   Joct �$  @I� �$  �K[)  �$   K�%  "�$   K�  &�$   KdO  )�$   K\=  ,�$   K�P  /�$    K�C  3�$   @IzS  6�$  �I�O  9�$  JK�?  <�$  I(  Q�%  �#  I�Q  V�%  IO  Y�%   H�9  i;#  Jin w�%  �%  Jout z�%   L;v  ��&  M�f&  G9�   G�  G�  G˭  G�  G^�  Gj  GL�  $Gڭ  G<�  "G3�  $ M�&  G��   G��  G��  Gʠ  G�  G٠  Gc�  G�m    Ў  �j   r  �j  N6�  �k  �u  k  q    �#  <�u  =�u  >�u  @qv  A|v  B�v  C�v  D�v  E�v  Fw  G!w  H6w  ks  4{'  O�{  7j'  G�p   Pdmy Pmdy Pymd Pydm  Qks  t'  ��    L�  HC(  R�k  K�'  GQ   G� Gʄ  Gih  G~  SSv  L�'  �O  LZw    MQ�'  G��   G+�  G�1    �  N�'  �'   ��  Y�j  AFv  ^��  �'  2(  q  q  q   Q�  <(  ��    ۝  �l(  T@�  ��j  ۝  e(  �    ד  ��(  ��  ��  � �k  �4  ��t  {�  k   U��  ��  B,  �   {'   H��  �B,  �A  ��w   ��  �u  Vid }  H�b  �q  H7# ��  9�q  � )  +)  �w  �   9�q  �<)  L)  �w  �w  �   9�q  �])  r)  �w  �-  �j  �   ,�{  �wz  �(  �)  �)  �w   ,]�  �L�  �(  �)  �)  �w   ,\�  ��  �!  �)  �)  �w   ,ń  %و  )  �)  �)  �w   ,&�  6ܫ  )  *  *  �w   ,�  G�  )  &*  ,*  �w   ,ڡ  W)�  �j  E*  K*  �w   ,v�  {ּ  �'  d*  j*  �w   ,e�  C�  �'  �*  �*  �w   We�  �(  �*  �*  �w  �j   XІ  ��}  �(  �(  �*  �*  �w   X�k  ��  �(  �(  �*  �*  �w   Xy  ��n  �!  �(  +  +  �w   X�  �;h  )  �(  @+  F+  �w   X�  �_�  )  �(  g+  m+  �w   Xz  ���  )  �(  �+  �+  �w   X�  ���  �j  �(  �+  �+  �w   X4n  ��  �'  	�(  �+  �+  �w   X"�  �!}  �'  
�(  ,  	,  �w   .�q  ��  ,  .,  �w  �-  �j   !T  q  Y�  �t    Z
�  Db�  �-  
�   Y�  d�j  �p  e�  q�  f�t  �{  gq  Z�  hq    i�j  �  j�  #�  k�j  ��  l�   �  m�j  $Ӎ  n�  (ס  o�j  ,s�  p�'  0b�  q�'  4گ  v�w  8}  x�t  Cҽ  z9-  D-  �w  �   [ѽ  �B,  Y-  d-  �w  �j   $[�  Ewo  w-  �-  �w  ]u   ,�  �i�  �w  �-  �-  �w  �w   9ҽ  ��-  �-  �w  �w   !T  q  Y�  �t    W�  1�w  �(  U�  ��  �1  �   {'   H��  ��1  �A  ��w   ��  �u  Vid }  H�b  �q  H7# ��  9�q  �c.  n.  �w  �   9�q  �.  �.  �w  �w  �   9�q  ��.  �.  �w  �-  �j  �   ,�{  �4�  8.  �.  �.  �w   ,]�  ��y  8.  �.  �.  �w   ,\�  �x  �!  /  /  �w   ,ń  %Qj  E.  +/  1/  �w   ,&�  6҅  E.  J/  P/  �w   ,�  G@~  E.  i/  o/  �w   ,ڡ  Wݑ  �j  �/  �/  �w   ,v�  {��  �'  �/  �/  �w   ,e�  ��  �'  �/  �/  �w   We�  �-  �/  �/  �w  �j   XІ  ��  8.  �-  0  0  �w   X�k  ��|  8.  �-  50  ;0  �w   Xy  ���  �!  �-  \0  b0  �w   X�  ��~  E.  �-  �0  �0  �w   X�  �+�  E.  �-  �0  �0  �w   Xz  �Ձ  E.  �-  �0  �0  �w   X�  �Ƥ  �j  �-  �0  �0  �w   X4n  ���  �'  	�-  1  %1  �w   X"�  �P�  �'  
�-  F1  L1  �w   .�q  Y�  a1  q1  �w  �-  �j   !T  q  Y�  �t   Z��  Db�  3  
�   Y�  d�j  �p  e�  q�  f�t  �{  gq  Z�  hq    i�j  �  j�  #�  k�j  ��  l�   �  m�j  $Ӎ  n�  (ס  o�j  ,s�  p�'  0b�  q�'  4گ  v�w  8}  x�t  Cҽ  z|2  �2  �w  �   [ѽ  ��1  �2  �2  �w  �j   $[�  E8�  �2  �2  �w  ]u   ,�  �~w  �w  �2  �2  �w  �w   9ҽ  ��2  3  �w  �w   !T  q  Y�  �t   �-  B,  �1  U�  ,�  �3  �(    ��  2u  9ѹ  5^3  n3  �w  �j  �   Wй  D(3  �3  �3  �w  �j   !T  q  Y�  �t    U��  ,�  4  �-    ��  2u  9ѹ  5�3  �3  �w  �j  �   Wй  D�3  �3  
4  �w  �j   !T  q  Y�  �t   U��  Z�  D6  �   Vid �}  H�b  `q  H�B  aD6  H7# b�  9��  pz4  �4  �w  �   -get �-�  O4  �4  �4  �w  O4  O4  �t  �u  �w  x   -get ��t  O4  �4  �4  �w  O4  O4  �t  �u  �w  	x   W��  �4  5   5  �w  �j   X�  l�z  D6  4  A5  e5  �w  O4  O4  �t  �u  �w  x   X�  yC�  D6  4  �5  �5  �w  O4  O4  �t  �u  �w  	x   /Ȋ  �_�  D6  �5  �5  Y�  �t  �w  O4  O4  �u  �w  �x   B4  /E�  �L�  D6  6  16  Y�  �t   �w  O4  O4  �u  �w  �x   !T  q  1�  D6   ��  2�7  !_   }'  C[_  (T  a_y   Fe  B8  �>  bo6  �b  @q  (� D�`  X�  f�6  �6  ey   X�  p�6  �6  ey  ky   X�  t�6  �6  ey  _y   /*  {p  �6  7  	7  qy   /�F  �C�  wy  !7  '7  ey   /�F  �ޙ  D6  ?7  J7  ey  �j   /|�  ���  �t  b7  m7  qy  }y   #  �%�  o6  �7  �7  qy   #��  Ú�  �t  �7  �7  qy   o6  !T  q  �E  !   4  U�  ��  �9  �   Vid |}  H�b  �q  H�B  ��9  H7# ��  90�   8  +8  x  �   -put ��  �7  D8  c8  x  �7  �t  �u  �7  st   -put 1��  �7  |8  �8  x  �7  �t  �u  �7  x   8  W/�  8�7  �8  �8  x  �j   X�  9i�  �9  �7  �8  9  x  �7  �t  �u  �7  st   X�  _:{  �9  �7  "9  A9  x  �7  �t  �u  �7  x   ,�  ���  �9  d9  ~9  Y�  �t  x  �7  �u  �7  x   �7  ,��  ���  �9  �9  �9  Y�  �t   x  �7  �u  �7  x   !T  q  1QJ  �9   ;G  �,;  �   }'  �[_  (T  �y   �U  �t  �E  ��`  "  �&:  1:  �y  �y   "  �A:  L:  �y  �y   /�  �'V  �y  d:  o:  �y  q   ,*  )A  �y  �:  �:  �y   ,�F  	j8  �y  �:  �:  �y  �j   ,�F  �8  �y  �:  �:  �y   ,V  �0  �t  �:  �:  �y   ,�E  L  �y  	;  ;  �y  �j  /M   !T  q  �E  !   �7  U�N  i�  �=  �   H��  r�=  \�A  u!x  Vid >}  H�b  oq  H7# p�  9��  ��;  �;  'x  �   9��  ��;  �;  'x  !x  �   9��  ��;  �;  'x  �-  �   ,�{  �w:  p;  <  <  -x   ,]�  ��H  p;   <  &<  -x   ,\�  �DU  �!  ?<  E<  -x   ,��  �  };  ^<  d<  -x   ,�p  �kV  };  }<  �<  -x   W�o  A1;  �<  �<  'x  �j   XІ  �n  p;  1;  �<  �<  -x   X�k  d�  p;  1;  �<  �<  -x   Xy  �  �!  1;  =  =  -x   X��  (��  };  1;  :=  @=  -x   X��  5P�  };  1;  a=  g=  -x   .��  E��  |=  �=  'x  �-   !T  q   Z0T  h �  �>  
�   Y�  "�j  �p  #�  q�  $�t  ��  %�j  ��  &�  �p  '�j  9i  (�   �{  )q  $Z�  *q  %3�  03x  &ݎ  6Cx  J}  8�t  d��  :T>  _>  Sx  �   [��  P�=  t>  >  Sx  �j   $[�  NC�  �>  �>  Sx  ]u   ,�  I��  Yx  �>  �>  Sx  _x   9��  L�>  �>  Sx  _x   !T  q   1;  �=  Ut�  R�  U?  1;   9��  Y?  *?  ex  �j  �   W��  h�>  @?  K?  ex  �j   !T  q   U�p  {�   G  �   Vid �}  H�b  �q  H�B  �D6  9mF ��?  �?  kx  �   -get ���  �?  �?  �?  qx  �?  �?  �u  �w  wx   -get �k�  �?   @  @  qx  �?  �?  �u  �w  }x   -get ��  �?  8@  W@  qx  �?  �?  �u  �w  �x   -get ���  �?  p@  �@  qx  �?  �?  �u  �w  �x   -get �B�  �?  �@  �@  qx  �?  �?  �u  �w  �x   -get ��  �?  �@  �@  qx  �?  �?  �u  �w  �x   -get �t�  �?  A  7A  qx  �?  �?  �u  �w  �x   -get y�  �?  PA  oA  qx  �?  �?  �u  �w  �x   -get �  �?  �A  �A  qx  �?  �?  �u  �w  �x   -get S�  �?  �A  �A  qx  �?  �?  �u  �w  x   -get 6݋  �?  �A  B  qx  �?  �?  �u  �w  �x   WK�  <U?  -B  8B  kx  �j   /R�  �Դ  D6  PB  oB  qx  D6  D6  �u  �w  �x   X�  M��  D6  U?  �B  �B  qx  �?  �?  �u  �w  wx   X�  �q�  �?  U?  �B  �B  qx  �?  �?  �u  �w  }x   X�  �G�  �?  U?  C  /C  qx  �?  �?  �u  �w  �x   X�  ��  �?  U?  PC  oC  qx  �?  �?  �u  �w  �x   X�  ���  �?  U?  �C  �C  qx  �?  �?  �u  �w  �x   X�  ���  �?  U?  �C  �C  qx  �?  �?  �u  �w  �x   X�  �%�  �?  U?  D  /D  qx  �?  �?  �u  �w  �x   X�  ���  D6  	U?  PD  oD  qx  �?  �?  �u  �w  �x   X�  ��  D6  
U?  �D  �D  qx  �?  �?  �u  �w  �x   X�  �p�  D6  U?  �D  �D  qx  �?  �?  �u  �w  x   X�  ��  D6  U?  E  /E  qx  �?  �?  �u  �w  �x   ]�f  Is  ME  bE  |�  q  qx  �j  �  q   y?  ,�e  q��  D6  �E  �E  ]T  %   qx  D6  D6  �u  �w  }x   ,f�  q��  D6  �E  �E  ]T  �j  qx  D6  D6  �u  �w  �x   ,��  qF�  D6  F  *F  ]T  k  qx  D6  D6  �u  �w  �x   ,�  q^�  D6  LF  kF  ]T  7   qx  D6  D6  �u  �w  �x   ,�h  q�  D6  �F  �F  ]T  0k  qx  D6  D6  �u  �w  �x   ,��  qº  D6  �F  �F  ]T  )k  qx  D6  D6  �u  �w  �x   !T  q  1�  D6   U?  U"(  ��  *M  �   Vid �	}  H�b  �q  H�B  ��9  9H �TG  _G  �x  �   -put �F!  6G  xG  �G  �x  6G  �u  )G  �t   -put 	&"  6G  �G  �G  �x  6G  �u  )G  %    -put #	z"  6G  �G  �G  �x  6G  �u  )G  7    -put )	�"  6G  H  +H  �x  6G  �u  )G  0k   -put -	;#  6G  DH  ^H  �x  6G  �u  )G  )k   -put ^	�!  6G  wH  �H  �x  6G  �u  )G  zt   -put b	/K  6G  �H  �H  �x  6G  �u  )G  st   -put w	=I  6G  �H  �H  �x  6G  �u  )G  l   .&�  ���  I  5I  �x  �j  �  q  �j  k  k  �x   .V�  A{|  JI  sI  �x  �j  �  q  �u  k  k  �x   .å  �  �I  �I  �x  q  /M  �u  k  �j  �x   W�  �	G  �I  �I  �x  �j   X�  @5�  �9  G  �I  J  �x  6G  �u  )G  �t   X�  �	�s  6G  G  )J  CJ  �x  6G  �u  )G  %    X�  �	��  6G  G  dJ  ~J  �x  6G  �u  )G  7    X�  �	>�  6G  G  �J  �J  �x  6G  �u  )G  0k   X�  �	�f  6G  G  �J  �J  �x  6G  �u  )G  )k   X�  t��  �9  G  K  /K  �x  6G  �u  )G  zt   X�  ���  �9  G  PK  jK  �x  6G  �u  )G  st   X�  ���  �9  	G  �K  �K  �x  6G  �u  )G  l   ,	�  M�  �9  �K  �K  ]T  %   �x  �9  �u  q  %    ,�  Mf  �9  L  L  ]T  7   �x  �9  �u  q  7    ,��  M�  �9  ?L  YL  ]T  0k  �x  �9  �u  q  0k   ,3�  M6�  �9  {L  �L  ]T  )k  �x  �9  �u  q  )k   ,�  ���  �9  �L  �L  ]T  zt  �x  �9  �u  q  q  zt   ,��  ��  �9  �L  M  ]T  st  �x  �9  �u  q  q  st   !T  q  1QJ  �9   G  �>  b�  ^��  ��  �O  �   ��  ��O  _�A  ��x  _`|  ��-  _^�  ��j  Vid B}  +�  ��M  �M  �x  �   +�  ��M  �M  �x  �x  �   +�  ��M  �M  �x  �-  �j  �   .�E  Ke�  N  N  �x  k  �  �j  �v   `��  �c�  3N  >N  �x  �x   `��  �?�  RN  ]N  �x  �x   `�  �j  qN  |N  �x  �x   `k�  ���  �N  �N  �x  �j   `ѭ  ��  �N  �N  �x  �x   `��  �v  �N  �N  �x  �x   .��  П  �N  �N  �x  �x   .��  ��  O  O  �x  �x   .*�  (L�  .O  9O  �x  �x   W�  ::M  OO  ZO  �x  �j   .ƙ  G��  oO  zO  �x  �-   !T  q   a�  �;�  �R  
�   !�  ��x  ��  @�j  w�  A�j  �m  B�j  ��  C�j  �  D�j  @�  E�j  ��  F�j   ^�  G�j  $k�  H�j  (7�  K�j  ,*l  L�j  0l�  M�j  4�l  N�j  8�v  O�j  <͋  P�j  @Ջ  Q�j  D�  T�j  H�  U�j  Lε  V�j  PR�  W�j  Tb�  X�j  X[�  Y�j  \��  Z�j  `=q  ]�j  d�  ^�j  hHq  _�j  l�  `�j  pSq  a�j  t^q  b�j  xiq  c�j  |tq  d�j  �q  e�j  ��  f�j  �s  g�j  �y�  h�j  �n�  k�j  ���  l�j  ���  m�j  �ۻ  n�j  ���  o�j  �Ɂ  p�j  ���  q�j  ��  r�j  ��  s�j  �ͮ  t�j  �{�  u�j  ���  v�j  �}  x�t  �b�  z�Q  �Q  �x  �   c�  ��O  R  R  �x  �j   $[�  ��f  1R  <R  �x  ]u   /�  ���  �x  TR  _R  �x  �x   +�  �oR  zR  �x  �x   !T  q   :M  �O  U|  ��  �S  �   Vid '}  H�b  �q  H�B  ��9  9�p  ��R  �R  y  �   -put v��  �9  S  %S  y  �R  �u  �R  �v  �j  �j   -put �x  �R  >S  bS  y  �R  �u  �R  �v  q  q   W�p  �R  xS  �S  y  �j   X�  �ي  �9  �R  �S  �S  y  �R  �u  �R  �v  q  q   !T  q  1QJ  �9   �R  U�n  +�  MT  �R   9^�  3	T  T  y  �j  �   W]�  9�S  /T  :T  y  �j   !T  q  1QJ  �9   UC�  p�  �X  �   2'   Vid �}  H�b  vq  H�B  wD6  9��  ��T  �T  y  �   ,ݚ  ���  >'  �T  �T  y   ,g�  �x  �T  �T  U  y  �T  �T  �u  �w  �v   ,C�  �N�  �T  U  =U  y  �T  �T  �u  �w  �v   ,�  ���  �T  VU  uU  y  �T  �T  �u  �w  �v   ,�  d  �T  �U  �U  y  �T  �T  �u  �w  �v   ,��  s�  �T  �U  �U  y  �T  �T  �u  �w  �v   W��  "MT  �U  V  y  �j   Xښ  l��  >'  MT  'V  -V  y   Xd�  3g  D6  MT  NV  mV  y  �T  �T  �u  �w  �v   X@�  
�  D6  MT  �V  �V  y  �T  �T  �u  �w  �v   X�  '�  D6  MT  �V  �V  y  �T  �T  �u  �w  �v   X	�  C5t  D6  MT  W  -W  y  �T  �T  �u  �w  �v   X��  _��  D6  MT  NW  mW  y  �T  �T  �u  �w  �v   , t  I��  D6  �W  �W  y  �T  �T  �x  �j  �j  �  �u  �w   ,r  t׵  D6  �W  �W  y  �T  �T  �x  �x  �  �u  �w   ,m}  �,y  D6  X  8X  y  �T  �T  �x  �x  �  �u  �w   ,��  s>�  D6  QX  uX  y  �T  �T  �u  �w  �v  �j   xT  !T  q  1�  D6   MT  U��  ��  �X  MT   9Z�  ��X  �X  #y  �j  �   WY�  ��X  �X  �X  #y  �j   !T  q  1�  D6   Ul�  ��  K[  �   C(   \l�  ��-  \��  ��j  Vid H}  H7# ��  9�@  �dY  oY  )y  �   9�@  ��Y  �Y  )y  �-  �j  �   ,@�  ���  P(  �Y  �Y  /y  $u  ]u   ,@�  ���  P(  �Y  �Y  /y  $u  ]u  �j   -get ���  FY  Z  Z  /y  P(  �j  �j  5y   FY  .<_  ޏ  9Z  DZ  /y  P(   W�  �X  ZZ  eZ  )y  �j   X=�  eu  P(  �X  �Z  �Z  /y  $u  ]u   X�  MUo  �!  �X  �Z  �Z  /y  P(  �j  �j  ;y   d`�  4
h  �X  �Z  �Z  /y  P(   ,(h  8_�  k  [  [  /y  5y   ,�  @ck  FY  6[  A[  /y  k   !T  q   �X  �!  Um�  W�  �[  �X   +�f  P}[  �[  Ay  �j  �   W�f  bU[  �[  �[  Ay  �j   !T  q   U~�  ��  .\  .\   9��  ��[  �[  Gy  �j  �   W��  ��[  \  \  Gy  �j   3�  q  �e  q  �$  �l   8(�  D\  Vid a}   U_}  H�  i^  �   \�t  U�-  Vid �}  H7# O�  93  c�\  �\  My  �   93  q�\  �\  My  �-  �   ,��  ��  �j  �\  �\  Sy  �j  �j  �j  �j   ,~  �n�  v\  ]  ]  Sy  �j  �j   ,#�  ���  %   5]  E]  Sy  �j  �j   ,��  ���  �j  ^]  n]  Sy  �j  �j   , ~  ���  �  �]  �]  Sy  k  �j  �   W�  �D\  �]  �]  My  �j   X	�  ��  �j  D\  �]  �]  Sy  �j  �j  �j  �j   X*k  �?�  v\  D\  ^  )^  Sy  �j  �j   X �  ��  %   D\  J^  Z^  Sy  �j  �j   v\  !T  q   D\  U��  ��  �^  D\   9�t   �^  �^  Yy  �j  �   W�t  n^  �^  �^  Yy  �j   !T  q   �  X!_  :	|  ���  _  �u  q  k  �j  /M  /M   !T  q  �E  !   ��  v[_  �#  �  e_Tp q  �.  0k  �?  k  �   �t   8�M  �`  ,�* �e  �z  }_  �_  �z   �b  �q  ,�* �_e  �z  �_  �_  �z   .cb  �Pc  �_  �_  {  �j   ,�-  �  �z  �_  �_  �z   ,�-  P  �z  `  `  �z   .� !4  !`  ,`  {  �j   ,�c  <�c  K`  E`  K`  {   Fe  �8  ,�a  R(b  K`  p`  v`  {   ,�S  �YH  K`  �`  �`  {  �_   ,�W  �B  /M  �`  �`  {  ��  /M   �_  !T  q  1�E  !   2�Y  D6  2�8  �9  ��  ('a  #V�  +W�  �y  a  a  �y  ]u   f  �1   �`  ~  (da  #V�  +��  �y  Oa  Za  �y  ]u   f  B,   ,a  {  2�a  #V�  5��  �y  �a  �a  �y  ]u   f  �=   ia  �k  ��a  �q  ��  ��  ��  � ��j  �4  ��t  {�  �j   [_  f�*  �t#  b  t#  t#   8�+  �c  ,��  a�)  4b  )b  4b  ށ  q   H�b  �q  gis 1�c  �t  Xb  hb  ށ  "  q   //�  �^�  �j  �b  �b  ށ  "  �j  �j   ,g�  ��  q  �b  �b  ށ  4b  q   ,k�  ��  4b  �b  �b  ށ  4b   XKC  3�T  4b  b  c  c  ށ  q   X҉  d�  q  b  /c  ?c  ށ  4b  q   XKC  J��  �j  b  `c  uc  ށ  �j  �j  �   ,��  |�  �j  �c  �c  ށ  �j  �j  �   Vid �}  7+3  ��3  �c  ށ    b  �  f*  K�"  �c  �"  �"   ff3  p�9  d  !T  q  �9  �j  �j   f��  ҧt  >d  !T  q  �E  !  }y  }y   f	W  ��  Xd  �  t#   t#  fͳ   �<�  �d  e_Tp 7   <�  <�   f l  ̧t  �d  !T  q  �E  !  }y  }y   f�*  O�"  �d  �"  �"   f+  W�"  �d  �"   f}�  ��t  �d  e_Tp q  �t  �t   f�  ɲa  e  8�  �j  �y   fz�  !Z�a  De  ��  �j  �j  �j  �   f|�  !r�a  ge  f�  �j  �j  �j   0��  8��  �j  �e  |�  k  �j  �j  h �-  0}`  ��d  l�  �e  �R  b  ]u   0�  ��u  |�  �e  �R  .\  ]u   .\  09p  ���  �   f  �R  D\  ]u   0�~  ��j  ��  "f  �R  1;  ]u   0��  �Ҁ  ��  Df  �R  G  ]u   0c�  ��w  <�  ff  �R  U?  ]u   0:�  ���  ��  �f  �R  �-  ]u   0�v  �ٮ  t �f  �R  �(  ]u   0=�  ��h  % �f  �R  �7  ]u   0�  �F�  � �f  �R  4  ]u   0�  �Ü  3 g  �R  :M  ]u   0h�  ��  3 2g  �R  �R  ]u   0r�  �H�  � Tg  �R  MT  ]u   0�  ��  A vg  �R  �X  ]u   0/�  h��  �t  �g  �R  b  ]u   0α  h/�  �t  �g  �R  .\  ]u   0��  hϞ  �t  �g  �R  D\  ]u   0w�  h��  �t  �g  �R  1;  ]u   0�g  hL�  �t   h  �R  G  ]u   09�  h|�  �t  Bh  �R  U?  ]u   0��  h�v  �t  dh  �R  �(  ]u   0�m  h2l  �t  �h  �R  �7  ]u   0ڌ  hz  �t  �h  �R  4  ]u   0zj  h�g  �t  �h  �R  :M  ]u   0�r  h�{  �t  �h  �R  �R  ]u   0,�  h�~  �t  i  �R  MT  ]u   0�  hþ  �t  0i  �R  �X  ]u   Jm  ���  k  li  !T  q  k  q  �j  �  �j  �j   @w  s�  �j  �i  !T  q  ]T  7   k  7   �j  �#  �t   /M  !�  q�  �j  �i  !T  q  ]T  )k  k  )k  �j  �#  �t   i	@  "8�N  ��  "N)�  j  �j  h 0��  �Ki  �t  5j  �j  �  ;y   �  R�l  Yj  �j  x  �w  |�   h�  H!o  }j  �j  �x  �w  |�   j<�  M��  �j  �x  �w  |�    f)%  Kk  �j  �j  �j   kint �j  q  lGT  P�j  >   m�p  q  �  #�j  �  �  o  �	  �  qW  #!�j    #")k  �  #  .  $<k  `  $D�j  �  $Wk  �  $_k  �  $e�j  t   $m�j  a  $u�j    $~�j  �  $��j  3  $��j  �  $��j  H  $��j  y  $��j    $��j  s  $��j  T   $ȸj  �  $иj  F  $׸j  �  $�j  �  $�j    $�j  V  $�j  �  ns  %N�j  �  %V�j  \	  &2�j  o  &7�j  �  &<�j  �  &C�j  �  '�j  �l  op(pO qO (!�l  q$   Est  Ų  )Y�l  |  )Z7    ��  )]�l  |  )^)k   �  +$,,�  ,-�  K  ,:zn  �e  ,=�  � ,?k  "  ,@�j  �4  ,A�t  �J  ,B�t  �A  ,OAm  Gm  �t   �A  ,QWm  bm  �t  �t   �A  ,Vrm  }m  �t  �j   /�
 ,Y51  m  �m  �m  �t  m   /�
 ,]�R  m  �m  �m  �t  %m   /� ,c?  m  �m  �m  �t  �l  l   `_ ,m.   �m  n  �t  m  �l   /�3  ,q89  �l  'n  -n  �t   `.E  ,��3  An  Qn  �t  m  �t   `�(  ,��(  en  pn  �t  m   e_Tp q   �l  LZD  -��p  \F�  -�k   H��  -�x(  H�4  -��(  H� -��(  *��  -��n  �n  jw   9��  -��n  �n  jw  pw   ,*  -��}  �n  o  o  {w   ,Ư  -�?s  �n  ,o  2o  {w   ,�F  -�Ϭ  �w  Ko  Qo  jw   ,�F  -��  n  jo  uo  jw  �j   ,a�  -�
�  �w  �o  �o  jw   ,a�  - ��  n  �o  �o  jw  �j   ,�:  -,�  �n  �o  �o  {w  �n   ,�F  -		n  �w  �o   p  jw  �n   ,(*  -��  n  p  $p  {w  �n   , I  -h�  �w  =p  Hp  jw  �n   ,�O  -7k  n  ap  lp  {w  �n   ,WC  -]�  pw  �p  �p  {w   {�  k  �  �   L8E  -��r  \F�  -��j   H��  -��a  H�4  -��a  H� -��a  *��  -��p  �p  �y   9��  -�q  q  �y  �y   ,*  -���  �p  ,q  2q  �y   ,Ư  -�p�  �p  Kq  Qq  �y   ,�F  -�5�  �y  jq  pq  �y   ,�F  -�÷  �p  �q  �q  �y  �j   ,a�  -��j  �y  �q  �q  �y   ,a�  - �i  �p  �q  �q  �y  �j   ,�:  -m�  �p  �q  �q  �y  �p   ,�F  -	�u  �y  r  r  �y  �p   ,(*  -�  �p  8r  Cr  �y  �p   , I  -*�  �y  \r  gr  �y  �p   ,�O  -�  �p  �r  �r  �y  �p   ,WC  -�i  �y  �r  �r  �y   {�  �j  �  �   �q  )5�r  |  )67   YX�  �t  H�  7   ��  )k   n  s  )/s  |  )0�j   k�  )/&s  |  )0�j   h�  )?Gs  |  )Es  e_Tp �j   �}  )/_s  |  )0k   �  )?�s  |  )ESs  e_Tp k   k  )/�s  |  )07    sh  )?�s  |  )E�s  e_Tp 7    �  )/�s  |  )0)k   ��  )?�s  |  )E�s  e_Tp )k   �p  rU  
A�t  t  �y  �j   r9+  
N�t  +t  �y  �j   s�y  -��n  Xt  {�  k  �  �  ��  ��   t��  )��t  �  �j  �j    �� �� �� q2*  *7�t  u*8�   v-  v]  �  ]  -  v�  vq  v�j  �l  vzn  zn  �  v    �  . �j  �j  �t  �  �  �  �  v�  v�  v�  w7   ;u  x �  _  Lu  Ru  �j  �  v�!  �!  }  v�!  �!  �u  �!  k  wuu  �u  x w�u  �u  x �u  uu  v�!  �!  7   v�#  v�&  �l  /%   j�  /#%   ytm ,/,qv  ,g  /.�j   �  //�j  �  /0�j  ��  /1�j  ��  /2�j  ��  /3�j  ��  /4�j  �  /5�j  d�  /6�j   ��  /7%   $~�  /8�j  ( l\�  />�u  fѯ  /Hzt  �v  �u  �u   f��  /M�u  �v  �v   �u  f�  /C�u  �v  �v   �u  f#�  /ak  �v  �v   �v  �u  f�� /fk  w  w   w  �u  f��  /W�v  !w  w   f[v  /\�v  6w  w   f��  /R,   Zw  k  ,   �j  �v   wq  jw  z)l   n  vvw  k  �r  vn  �(  �(  �j  �-  .  �-  3  wq  �w  z)l  
 B,  vB,  v3  �1  v�1  v#3  (3  �3  4  �7  v�#  vst  v\4  �7  ,;  v�8  I;  1;  �>  wq  Cx  z)l  # wq  Sx  z)l   �=  v�=  v�>  �>  U?   G  v�t  v%   v�j  vk  v7   v0k  v)k  v�t  vzt  v0l  v�!  G  *M  v�j  QM  :M  �R  �j  w�j  �x  z)l   �O  v�O  v�R  �R  �S  �S  MT  �X  �X  �X  K[  vZ  vP[  U[  �[  D\  i^  n^  W6  D6  v�6  �`  vD6  v�`  �9  �9  v
:  v�9  �`  #3  'a  3  da  �>  �a  %   �p  vRu  �s  v�p  �t  {�s  z  |XF  
A�y  |\;  
A�j  }~�T  
C�t    I  $z  /z  �h  /z   u  �  Bz  Mz  �h  /z   r  [z  fz  �h  /z     tz  z  �h  z   u  �  �z  �z  �h  �z   ;u  {�  �z  }�__p 	�0l    �  �z  �z  �h  �z   �_  �a  d_  �z  �z  �h  �z   �z  �_  {  {  �h  �z   [_  �_  +{  C{  �h  C{  �__n ��j   {  �_  V{  a{  �h  �z   �_  o{  z{  �h  �z   `  �{  �{  �h  C{  �__n !�j   *  �{  �{  �h  z   n3  �{  �{  �h  �{  �#  �t   �w  �3  �{  |  �h  |  �#  �t   �w  �4  |  ,|  �h  ,|  �#  �t   �w  �8  ?|  T|  �h  T|  �#  �t   x  *?  g|  ||  �h  ||  �#  �t   ex  B  �|  �|  �h  �|  �#  �t   kx  �I  �|  �|  �h  �|  �#  �t   �x  bS  �|  �|  �h  �|  �#  �t   y  T  }  }  �h  }  �#  �t   y  �U  /}  D}  �h  D}  �#  �t   y  �X  W}  l}  �h  l}  �#  �t   #y  {t  �}  |XF  
N�y  |\;  
N�j   �  �}  �}  �h  z  �__a 	�}   �t  �[  �}  �}  �h  �}  �#  �t   Ay  �^  �}  ~  �h  ~  �#  �t   Yy  �  ~  %~  �h  %~   u  O  8~  l~  �h  /z  �%  	S�  �Q  	S�  }��c  	Uu    �  z~  �~  �h  /z  �%  	A�  �__s 	A�j   �[  �~  �~  �h  �~  �#  �t   Gy  {C  �~  |hR  ��~  |mR  ��~   �t  �t  a       �h  z   C    0  �h  z  �__n 	��     >  I  �h  /z   {�  {  �__s 
�t  �__n 
�  �__a 
{   �t  {"  �  ��e  �t  ��e  �t  �__n �   {�  �  �__d 	dk  �__s 	d�j  �__n 	d�   {j  �  �__c �   �t  {�  �  �__c  �   �t  ,`  ,�  F�  �h  C{  }��&  >K`    W`  T�  n�  �h  C{  }��&  TK`    v`  |�  ��  �h  C{  �__c ��_  }��&  �K`    {�  Ȁ  �hR  $Ȁ  �mR  $̀   �t  �t  �  ��  �  �h  �   iu  {�a  �  �__a �t#  �__b �t#   �&  �#  '�  2�  �h  2�   �  �#  �#  K�  r�  �h  r�  ��%  2�#  }�'U  4�#    7�  $  ��  ��  �h  2�   %$  ��  ��  �h  2�   D$  ��  ށ  �h  r�  ��R  �/M  }�'U  �/M    �c  b  �  
�  �h  
�  �__c aq   ށ  Ab  �  }�  �h  
�  �__m 2"  �__c 2q  }~�&  8�t  ~�`  9�c  ~�b  :�  }~a  =+"  }~�c  @�t      hb  ��  ��  �h  
�  �__m �"  |�a  ��j  |�a  ��j   �  �  ̂  �  �h  �  �4&  r�   ��  �R  ��  �  �h  �|  �4&  ��   a  �  (�  �h  /z   {�c  K�  �__a K�"  �__b K�"   {F  }�  �__s �t  �__n �  �__a -   h$  ��  ��  �h  2�   {'  �2(  H��  ��  �h  ��   ��  2'  �j'  4Ճ  ��  �h  ��   ��  �T  �  �  �h  D}  �4&  ��   C(  �\(  �#�  .�  �h  .�   �  ��  /E  Q�  ��  |�  q  �h  ��  �j  �R'  I�  �__c Iq  }��&  K�j    qx  �b  ��  ф  �h  
�  �__c �4b  ��  �q  }�__t ��j    o:  ߄  �  �h  �   �y  �:  ��  �  �h  �   1m  �  !�  �h  !�   �t  6  4�  ?�  �h  ?�   �t  bm  R�  g�  �h  !�  �#  �t   g  u�  ��  �h  ?�  �#  �t   �n  ��  ��  �h  ��  �__i -���   jw  pw  �`  �`  ΅  �  �h  C{  �__s ���  �__n �/M   {�  �  �__s �t   {�c  A�  !T  q  �__s p�9  |�+  p�j  |R'  p�j   �7  O�  g�  �h  g�  }~�^  ŧ7    qy  �6  z�  ��  �h  g�   	7  ��  ��  �h  ��   ey  {d  ؆  !T  q  �E  !  �__a �؆  �__b �݆   }y  }y  vXd  vt#  {>d  �  �__a ��  �__b �t#   �  �b  $�  <�  �h  
�  �__c 4b   v�u  {]d  n�  e_Tp 7   �__a  �n�  �__b  �s�   <�  <�  �N  ��  ��  �h  ��  �b�  �x   �x  �N  ��  Ǉ  �h  ��  |b�  ��x   ]N  Շ  �  �h  ��  ||�  ��x   N  ��  �  �h  ��  |q~  ��x   >N  �  3�  �h  ��  |�  ��x   {�d  h�  !T  q  �E  !  �__a �h�  �__b �m�   }y  }y  lp  ��  ��  �h  ��   {w  �  ��  ��  �h  /z   v�r  {+t  �  {�  k  �  �  �\C  -��  �?)  -��   ��  ��  Gm  ��  �  �h  !�  �   �t  L  !�  8�  �h  ?�  �__a s8�   �t  �  K�  V�  �h  /z   ��  	h�  }�  �h  }�  �#  �t   u  r)  ��  ��  �h  ��   �w  �)  ��  ��  �h  ��   ,*  ǉ  ҉  �h  ��   �)  ��  �  �h  ��   �
  ��  �  �h  %~  �#  �t   �)  �  '�  �h  ��   �)  5�  @�  �h  ��   *  N�  Y�  �h  ��   K*  g�  r�  �h  ��   j*  ��  ��  �h  ��   �.  ��  ��  �h  ��   �w  �.  ��    �h  ��   o/  Њ  ۊ  �h  ��   �.  �  �  �h  ��   /  �  �  �h  ��   1/  �  &�  �h  ��   P/  4�  ?�  �h  ��   �/  M�  X�  �h  ��   �/  f�  q�  �h  ��   &<  �  ��  �h  ��   -x  E<  ��  ��  �h  ��   d<  ��  ��  �h  ��   �;  ϋ  ڋ  �h  ��   <  �  �  �h  ��   D>  �  �  �h  �  �4&  :�   Sx  {�d  A�  �__a O�"  �__b O�"   {�d  X�  �__a W�"   �  f�  ��  �h  }�  �v�  	k  �__a 	��   �t  ��	  �	  ��  ��  �h  %~   c  ��  ֌  �h  %~  �__c 	�q   n  �  �  �h  /z   �  ��  �  �h  %~  �%  	U�   z  #�  .�  �h  %~   �  <�  T�  �h  %~  �__n 	��   �  b�  m�  �h  /z     {�  ��  �h  %~  �__n 	��  �__c 	�q     ��  ƍ  �h  %~  ��^  	�ƍ   $u  �$  ٍ  �  �h  2�   S  �  ��  �h  %~   {�d  �  e_Tp q  �   �   �t  �t  {�d  >�  8�  �j  >�   �y  {e  r�  ��  �j  |z  !Z�j  |�l  !Z�j  �   {Xt  ��  �  �j  |Ő  )��j   {De  ��  f�  �j  |z  !r�j  |�l  !r�j   {Z	  �  �__p 	�k  �۶  	��j  �nh  	��j   {�  A�  ß  �j  |�|  |�j  |�h  |�j  �__a |A�  �  }~�  ��  �__r �u    �t  {"  ��  �  �j  ��|  	��j  ��h  	��j  �__a 	���  �  � �t  {T  ʏ  �  �j  ��|  	��j  ��h  	��j  �__a 	�ʏ  � �t  �  �  �  f�  �j  �h  %~  |�|  �j  |�h  �j  �__a ��   �t  �  &�  1�  �h  /z   �^�  W�  �w  B�j  �-�  B�j   �b  e�  }�  �h  
�  �__c 3q   �W�  �T  ��   ���  ��  �e�  � �o�  � c  ��  ߐ  �h  
�  �__c d4b  ��  dq   ���  �  ��   ���  �  ���  � �Đ  ��ѐ  � �*  %�  0�  �h  ��   ��  �}  ��   �L�  V�  �%�  �  �*  d�  o�  �h  ��   �V�  �  ��   ���  ��  �d�  �  �+  ��  ��  �h  ��   ���  ��  ��   �ʑ  ԑ  ���  �  �+  �  �  �h  ��   �ԑ  �  ��   �	�  �  ��  � �+  !�  ,�  �h  ��   ��  !}  ��   �H�  R�  �!�  � �/  `�  k�  �h  ��   �R�  �  �   ���  ��  �`�  �  0  ��  ��  �h  ��   ���  �|   �   �ƒ  В  ���  �  �0  ޒ  �  �h  ��   �В  Ƥ  0�   ��  �  �ޒ  �  �0  �  (�  �h  ��   ��  ��  @�   �D�  N�  ��  � %1  \�  g�  �h  ��   �N�  P�  `�   ���  ��  �\�  � ��{  Ń  ��   ���  Ó  ��{  � ����� �   ��{  �l  ��   �ߓ  ��  ��{  � ����� �   �<  �  �  �h  ��   ���  �n  ��   �.�  8�  ��  �  �<  F�  Q�  �h  ��   �8�  d�  ��   �m�  w�  �F�  �  �Y|  �  ��   ���  ��  �g|  � ����� �   �V  ��   �Ŕ  Ӕ  �h  Ӕ  �  y  �eZ  @��   ��  �  �h  �  � ��  ���  � /y  $u  ]u  ��Z  K��   �;�  R�  �h  �  � �P(  � �)^  � �!   �l�  ��  �h  ��  � ��k  ��j  W�  �:�  ��j  ��  ��-  �\;  7   ��    Sy  �	|  ��  0�   �Օ  �  �|  � �?��� �   �1|  �  @�   ��  %�  �?|  � �O��� �   ��|  ��  P�   �A�  [�  ��|  � �_��� �   ��|  �  `�   �w�  ��  ��|  � �o��� �   �Q   ��  ��  �h  ��  �#  �t   �x  ���  ��  p�   �Ֆ  �  ���  � ���� �   ��|  :�  ��   ��  %�  ��|  � ����� �   ��|  ��  ��   �A�  v�  �}  � ��|  ��   9��|  � ����� �    �!}  <�  ��   ���  ��  �/}  � ����� �   �I}  ��  ��   �ȗ  ��  �W}  � �!}  ��   ��/}  � ����� �    �*  �  �  �h  ��   ���  �n  ��&   �2�  B�  ��  ���� +  P�  [�  �h  ��   �B�  ;h  ��&   �w�  ��  �P�  ��� F+  ��  ��  �h  ��   ���  _�   �&   ���  ̘  ���  ��=� m+  ژ  �  �h  ��   �̘  ��  P�&   ��  �  �ژ  ��m� ;0  �  *�  �h  ��   ��  ��  ��&   �F�  V�  ��  ���� b0  d�  o�  �h  ��   �V�  �~  ��&   ���  ��  �d�  ���� �0  ��  ��  �h  ��   ���  +�  ��&   �Й  ��  ���  ���� �0  �  ��  �h  ��   ���  Ձ  �&   ��  %�  ��  ��-� �<  3�  >�  �h  ��   �%�  �  @�&   �Z�  j�  �3�  ��]� =  x�  ��  �h  ��   �j�  ��  p�&   ���  ��  �x�  ���� @=  ��  Ț  �h  ��   ���  P�  ��&   ��  ��  ���  ���� D-   �  �  �h  �  �#  �t   �w  ���  Xp  ��m   �8�  p�  ��  � ����d ���d ���d �-��d �=� �2   ~�  ��  �h  ��  �#  �t   �w  �p�  8�  @�m   ���  �  �~�  � �d��d �w��d ����d ����d ��� _>   ��  �  �h  �  �#  �t   ��  :�  ��Z   �+�  Y�  ���  � ����d ����d ����d �
� ���  �  �   �u�  ��  ��  � ���+�e  �p�  ,r  0�   ���  Ŝ  �~�  � �>��K�e  ��{  X�  P�!   ��  �  ��{  � ��{  X�   D�  ��{  �  �d� �q�e  ��{  M�  ��!   �7�  q�  ��{  � ��{  ��   Df�  ��{  �  ��� ���e  �	|  �s  ��!   ���  ǝ  �|  � �	|  ��   ���  �|  !�  ��� ���e  �1|  ki  ��!   ��  �  �?|  � �1|  ��   8�  �?|  @�  ��� ��e  ��  ��  �   �9�  S�  ���  � ���+�e  �Y|  ��  0�!   �o�  ��  �g|  � �Y|  8�   h��  �g|  _�  �D� �Q�e  ��|  8�  `�!   �Ş  ��  ��|  � ��|  h�   <��  ��|  ~�  �t� ���e  ��|  _m  ��!   ��  U�  ��|  � ��|  ��   �	J�  ��|  ��  ��� ���e  ���  6�  ��   �q�  ��  ���  � ������e  ��|  �  ��!   ���  �  ��|  � ��|  ��   ֟  ��|  ��  ��� ��e  ��|  e�  �!   ���  S�  �}  � ��|  �   9H�  �}  ۋ  ��|  �   9��|  ۋ  �$�  �1�e  �!}  m�  @�!   �o�  ��  �/}  � �!}  H�   "��  �/}  ��  �T� �a�e  �I}  ��  p�!   �Š  �  �W}  � �I}  x�   ��  �W}  �  �!}  x�   ��/}  �  ���  ���e  4b  ?c  /�  a�  �h  
�  ��k  J�j  �:�  J�j  �"y  J�   �!�  ��  ��"   �}�  ��  �/�  � �9�  ��F�  ��S�  ����#e  �DZ  ; ��  ҡ  �h  ҡ  �#  �t   )y  ���  }p  ��>   ��  �  ���  � ���  �������Ge  ���  D�  �   �9�  S�  ���  � ���+�e  ��}  ф  0�   �o�  ��  ��}  � �?�ס  �� �   ��}  8�  @�!   ���  �  ��}  � ��}  H�   cܢ  ��}  8�  �T�ס   �a�e  �]  ��  
�  �h  
�  �#  �t   My  ��  �g  p�>   �+�  U�  ���  � ���  ���������Ge  �9O  S f�  {�  �h  {�  �#  �t   �x  �U�  ��  ��m   ���  ڣ  �f�  � ���"  ����d ���  �
�����Ge  �U�  ��   �   ���  �  �f�  � �.��;�e  ��~  <  @�   �,�  F�  ��~  � �O��� �   ��~  ��  P�!   �b�  ��  ��~  � ��~  X�   ���  ��~  W�  �d� �q�e  ��}  ��2   ���  ,�  ��}  v�  ��}  ��  �q}  ���-  	�!�  ��}  �{}  ��  ��y  ���-  
V��y  ��y  ��  ��-  �	z  ݌     ����   ��]  ���'  �F�  _�  �h  ��  � ���  ��j  ����  ��j  ����  ��j  ��k~  ��j  ���-  T�  ���  �Z^  ��  ���  �Z^  ��  �__p ��j  ۍ  �u�  ��j  �  �__q ��j  S�  ���  ��j  ��  �Ϗ  ��.  ���  ��  ֎  ���  O�  ���  o�  ��  �k)  ���  ��.  ���  ֎  ���  O�  ���  o�  �.  �F�  ��.  	��s�  ֎  �f�  O�  �Y�  o�  �.  ����       �Ϗ  ��(.  �k�  ��  ��  ���  ��  ���  �  ��  �{)  ���  ��(.  ���  ��  ���  ��  ���  �  �(.  �F�  ��(.  	��s�  ��  �f�  ��  �Y�  �  �(.  ����       �@.  �  �/t  ��t  0�  ��  "�	   ���  ���  Y�  �+�[e  ��  +�h.  �ק  ���  l�  �5�[e  ��E]   ��  L��.  �Y�  ���  �  �4z  L��.  	# �  �Bz  �   ��}  R��.  	#��}  ��  ��}  ɐ  �����  �Rug   ��  Y��.  �Ш  ���  �  �4z  Y��.  	#��  �Bz  �   ��}  _��.  	#��}  �  ��}  1�  �����  �Rug   ��  ��   ��  �k)  �4z  ��   	#�  �Bz  �k)   ��}  ��   	#��}  O�  ��}  |�  �����  �PuL<�Rug    ���Ge  ��  ��@   �w�  ��  ��  ��  ���  �  ����c   ��}  ��  0�>   ���  ��  ��}  � ��  8�/  �  ���  �  �J�  �[��f� �n�Ge  ��  ��  p�F   ��  l�  ���  � ��  x�(/  �W�  ���  ;�  ���  ������ ���e ���Ge  ��}  �  ��F   ���  ��  ��}  � ��}  ��@/  �  ��}  q�  ��  ��@/  ���  q�  ���  ������  ���e ��Ge  O  �  -�  �h  %~  �__c 	-q  }�R'  	/�    ��]  ���  �G�  |�  �h  ��  ���k  ��j  ��:�  ��j  ��X/  q�  ��&  �v\  � ��^  �Z^  ��  �__p Ͽj  �  �u�  пj  }�  �R'  ��  ؓ  �__c �k  K�  �Ϗ  ��/  ͕�  ��  ��  ���  �  ���  O�  ��  �\/  ���  ��/  ���  ��  ���  �  ���  O�  ��/  �F�  ��/  	��s�  ��  �f�  �  �Y�  O�  ��/  �5��       ���  %�   ��  ���  ��  �X�  %�   	��}�  �p�  ��  �f�  ��    �`��   ɮ  �/t  ��  ĕ  ��  ��   �'�  ���  �  ���[e  ���  ���/    ��  2�  ��  ��/  ��  F�  �Mz  ���/  	/��  �[z  �4z  ��   	��Bz  �z  ��   	-�$z     ��~  ��   	2ѭ  ��~  e�  ��~  }�   �4z  ��   	3�  �Bz  �z  ��   	-�$z    �  ��-   	3��  �#  ��  �  ��  ���"   �#  ��  �  Җ  ��{  �   	�g�  ��{   ��~  �   	װ�~  ��~  �     ���3    �m�n]  ����d ���se ���n]  ����   ��  )��/  �@�  ���   �  �4z  )��/  	#�  �Bz   �   ��}  ,��/  	#��}  �  ��}  T�  �M���  �Rug   ��  d�   ���  ���  ��  �4z  d�   	#~�  �Bz  ��   ��}  j�   	#��}  ʗ  ��}  ��  �y���  �PuH<�Rug   �y�   *�  ���  �4z  y�   	#�  �Bz   ��}  ~�   	#��}  �  ��}  G�  �����  �Rug   �P�se �)��d �d��e ����e ����d ����e ����e  ���Ge  v�e  �ge  ���   ���  ���  � �%  8k  ���a  9�t  Z�  �-  :�j  �h�0  �'U  <k  ��  �gw  =k  ��  �X}  F�j  Ø  ��&  L�t  ��  � �/   [�  �R'  @�c  /�  �)�[e �4�se �A�#e �O��j   ����j  ���e �d��e �p��j  �x��d   |�  uc  ��  Ա  �h  
�  ��k  |�j  �:�  |�j  �"y  |�   ���  �  ���   ��  )�  ���  � ���  ����  ��Ʊ  ����#e ����c   ��  �c   �(  �E�  !�  ��  � �'�  ��3�  ��80  ��  �3�  �'�  �80  �@�  B�  �K�  �V�  k�  �`0  �b�  ��  ��0  �n�  ��  ����e ����e �+��e �]�f �y�"f ���7f ���Lf ���af ��vf �9��f      )  /�  G�  �h  G�  �4&  ��   �w  �!�  d�  P�L   �h�  ��  �/�  � �9�  ����  Q��0  ���  �ւ  ?�  �̂  v�   ��	,  ������Ge  +)  ͳ  �  �h  G�  ���  ��w  �4&  ��   ���  m  ��K   ��  n�  �ͳ  � �׳  ���  ����  ���0  �S�  �ւ  ��  �̂  �   ���	,  ������Ge  L)  |�  ��  �h  G�  �(�  ��-  �__s ��j  �4&  ��   �n�  ��  ��N   �ʴ  3�  �|�  � ���  ����  ����  ����  ��1  ��  �ւ  �  �̂  P�   �!�	,  �6��>�Ge  ���  wz  @�"   �O�  v�  ���  ��  ��  Q�   ��%�  ��    ���  L�  p�"   ���  ��  ���  Ŝ  �V�  ��   ��d�  �    �҉  ��  ��S   �յ  �  ���  ����  ��   ��  �  ���  ��  و   �S   ��  I�  ��  ��B�  �   &�P�  #�  �-�  �'�  ܫ  `�S   �e�  ��  �5�  ����  y�   7���  B�  ���  �@�  �  ��S   ���  ٶ  �N�  ��̘  ��   H�ژ  a�  ���  ���  )�   �"   ���  �  �ǉ  ��  ���  1�   X���  ��    �Y�  ּ  P�H   �8�  ^�  �g�  ��ԑ  h�   |��  ��    �r�  C�  ��H   �z�  ��  ���  ���  ��   ��!�  ޝ    R.  ��  Ʒ  �h  Ʒ  �4&  ��   �w  ���  �  ��L   ��  >�  ���  � ���  ����  ��81  �#�  �ւ  ��  �̂  4�   ��L1  �4��<�Ge  n.  L�  q�  �h  Ʒ  ���  ��w  �4&  ��   �>�  ��  @�K   ���  �  �L�  � �V�  ��c�  ����  A�h1  �Ҹ  �ւ  j�  �̂  ��   �n�L1  ������Ge  �.  ��  -�  �h  Ʒ  �(�  ��-  �__s ��j  �4&  ��   ��  ��  ��N   �I�  ��  ���  � ��  ���  ���  ����  ���1  ���  �ւ  מ  �̂  �   ���L1  ������Ge  ���  4�  ��"   �ι  ��  ���  D�  �R�  ��   ��`�  o�    ���  �y  �"   ��  8�  ���  ��  ���  !�   ����  ��    �ۊ  �x  @�S   �T�  ��  ��  ���  Y�   ��    �m�  ��  Qj  ��S   ���  Ⱥ  ��  ��V�  ��   &�d�  �  ���  ��  ҅   �S   ��  �  ��  ����  �   7���   �  �-�  �&�  @~  `�S   �,�  X�  �4�  ����  y�   H��  �  ���  �  ݑ  ��"   �t�  ��  �Њ  >�  �В  ��   X�ޒ  i�    �?�  ��  ��H   ���  ݻ  �M�  ���  �   |��  }�    �X�  ��  @�H   ���  �  �f�  ��N�  X�   ��\�  ��    )-  -�  E�  �h  �  �4&  z�   ��  �  ���   �a�  ��  �-�  � �7�  ����  ���1  ��ւ  ��̂  �   l2  ��  ��  �h  ��  �4&  z�   ���  Ք   ��   �ڼ  �  ���  � ���  ����   ��1  ��ւ  ��̂  �   M3  �  S�  �h  �{  �__s 5�j  �4&  5�  }�Y�  ;�-    ��  b�  ���   �o�  @�  ��  � �)�  ��  �6�  ��!�  ��2  6�  �9�  �  �/�  6�  ���  ��H2  �޽  �ւ  �  �̂  6�   ���	,  �t� � �*   %�  �D�  �\�1�3  �?�	,  �G�   �c��k�Ge �|�Ge  �3  N�  ��  �h  |  �__s 5�j  �4&  5�  }�Y�  ;�-    �@�  �  ���   ���  o�  �N�  � �X�  ��  �e�  ����  ��p2  6�  ���  ��  ���  
�  ���  ���2  ��  �ւ  ��  �̂  
�   ���L1  �D� ���*   T�  �s�  �\��3  ��L1  ��   �3��;�Ge �L�Ge  i4  }�  ��  �h  ,|  �4&  p�   �o�  �  P�   ���  �  �}�  � ���  ����  P��2  p�ւ  ��̂  �   ��4  p�>   � �  n�  �h  n�  ��__s �O4  ���h  �O4  ����  ��t  ��$  �s�  ���*  �x�  � �#�  �}�  �$ �w  �u  �w  x  ��4  ��>   ���  �  �h  n�  ��__s �O4  ���h  �O4  ����  ��t  ��$  ��  ���*  ��  � �{�  ��  �$ �u  �w  	x  8  %�  =�  �h  T|  �4&  �   ��  P�  ��   �Y�  ��  �%�  � �/�  ����  ���2  �ւ  ��̂  �   �+8  �@   ���  �  �h  �  ��__s �7  ����  �t  ��$  �  ���O  �7  ��#�  st  � x  �u  �c8  P�8   �(�  ��  �h  �  ��__s 1�7  ����  1�t  ��$  1��  ���O  2�7  ��{�  2��  � �u  x  �;  ��  ��  �h  ��  �4&  ��   'x  ���  M�  ��J   ���  .�  ���  � ���  ����  ��3  ��  �ւ  c�  �̂  ��   ���g=  ������Ge  �;  <�  a�  �h  ��  ���  �!x  �4&  ��   �.�  �  ��I   �}�  ��  �<�  � �F�  ��S�  ����  ��83  ���  �ւ  Т  �̂  �   ��g=  �!��)�Ge  �;  ��  �  �h  ��  �(�  ��-  �4&  ��   ���  ��  0�K   �,�  ��  ���  � ���  ���  ����  1�h3  �q�  �ւ  =�  �̂  t�   �^�g=  �s��{�Ge  ���  w:  ��"   ���  ��  �ϋ  ��  ���  ��   ���  գ    �ڋ  �H  ��"   ���  �  ��  �  �8�  ��   ��F�  �    �q�  DU  ��S   �.�  Z�  ��  ��%�  ��   ��3�  (�  ��  ���    @�S   �v�  ��  ���  ��j�  Y�   ��x�  G�  �m�  ���  kV  ��S   ���  ��  ���  ����  ��   ����  f�  ���  ��  f�   �S   ��  =�  ��  � ��  ����   ��3  ?�ւ  ��̂  �   	?  K�  �  �h  ||  �__s Y�j  �4&  Y�  }�Y�  _�-    �=�  D�  `��   ���  l�  �K�  � �U�  ��  �b�  ����  a��3  Z�  ���  ��  ���   �  ���  a��3  �
�  �ւ  ��  �̂   �   ���g=  �!� ���'   Q�  �p�  �\���3  ���g=  ���   ����Ge �)�Ge  �?  z�  ��  �h  �|  �4&  ��   �l�  ��  0�   ���  ��  �z�  � ���  ����  0�4  ��ւ  ��̂  �   ��?  P�8   ���  [�  �h  ��  ��e  ��?  ���h  ��?  ��$  �[�  ���*  �`�  ��__v �e�  �  �u  �w  wx  �7A  ��8   ���  ��  �h  ��  ��e  �?  ���h  �?  ��$  ��  ���*  ��  ��__v ��  �  �u  �w  �x  �oA  ��8   ��  e�  �h  ��  ��e  �?  ���h  �?  ��$  e�  ���*  j�  ��__v o�  �  �u  �w  �x  ��A  �8   ���  ��  �h  ��  ��e  �?  ���h  �?  ��$  ��  ���*  ��  ��__v ��  �  �u  �w  x  ��A  P�8   ��  o�  �h  ��  ��e  6�?  ���h  6�?  ��$  6o�  ���*  7t�  ��__v 7y�  �  �u  �w  �x  CG  ��  ��  �h  �|  �4&  ��   �~�  �  ��   ���  ��  ���  � ���  ����  ��84  ��ւ  ��̂  �   �_G  ��4   ��  ]�  �h  ]�  ��__s �6G  ��$  �b�  ���O  �)G  ��__v ��t  � �x  �u  �^H  ��6   ��  ��  �h  ]�  ��__s ^	6G  ��$  ^	��  ���O  ^	)G  ��__v ^	zt  � �u  ��H  0�:   ���  8�  �h  ]�  ��__s b	6G  ��$  b	8�  ���O  b	)G  ��__v c	st  � �u  ��H  p�2   �U�  ��  �h  ]�  ��__s w	6G  ��$  w	��  ���O  w	)G  ��__v x	l  � �u  ��M  * ��  ��  �h  {�  |4&  ��   ���  %s  ��R   ���  K�  ���  � ���  ����  ��X4  +&�  �ւ  Y�  �̂  ��   ���"  ���ZO  �����Ge  ��M  2 \�  }�  �h  {�  |��  ��x  |4&  ��   �K�  ^r  �Q   ���  �  �\�  � �f�  ��q�  ����  ��4  3��  �ւ  ƥ  �̂  ��   �6�"  �D�ZO  �Y��a�Ge  ��M  : �  X�  �h  {�  |(�  ��-  �__s ӿj  |4&  ��  }~R'  @�c  ~Y�  Ak    ��  ��  p��   �t�  U�  ��  � ��  ��(�  ��4�  ����  q��4  <��  �ւ  3�  �̂  j�   ��4  ��  �@�  ��  �K�  ��  ���[e ���se ���#e  ���"  ����f ���ZO  ���e ����Ge �'��e �>��d �F��e  ��  c�  P�   �q�  ��  ���  � ��  � ��  ?�  p�   ���  ��  ��  � �'�  � �Ǉ  j  ��   ���  ��  �Շ  � �߇  � �|N  ��   ���  �  �h  ��  � ���  ��j  Ҧ   ��N  ��   �0�  M�  �h  ��  � ���  ��x  � ���  v  ��G   �i�  |�  ���  � ���  � �x�  П  0 G   ���  ��  ���  � ���  � �N  ��  ��  �h  ��  ��  �x   ���  ��  � �   ���   �  ���  � ���  � O  �  &�  �h  ��  ��  (�x   � �  L�  �   �B�  U�  ��  � ��  � �Q  c�  y�  �h  ��  |4&  z�   �U�  ː  ��  ���  ��  �c�  � �m�  ����  ��4  ��ւ  ��̂  �   ��  #�  P   ���  �  ���  � ��  ����  P5  ��ւ  ��̂  �   �%S  p>   �6�  ��  �h  ��  ��__s �R  ��$  ��  ���O  �R  ��y  �v  ���l  q  ��!�  q  �  y  �u  �S  ��  ��  �h  }  �j  �4&  3�   ���  �o  �   ���  Y�  ���  � ���  ����  ���  �05  4��  ����  � ���  �05  ��ւ  ��̂  �    ��  p�  �   �u�  ��  ��  � ���  ����  �P5  ��ւ  ��̂  �   ��T  �   ���  ��  �h  Ӕ  � ���� �   ��T   8   ���  X�  �h  Ӕ  ���|  ��T  ���h  ��T  ��$  �X�  ���*  �]�  ��y  ��v  �  �u  �w  �U  @8   �z�  ��  �h  Ӕ  ���|  ��T  ���h  ��T  ��$  ���  ���*  ���  ��y  ��v  �  �u  �w  �=U  �8   ���  X�  �h  Ӕ  ���|  ��T  ���h  ��T  ��$  �X�  ���*  �]�  ��y  ��v  �  �u  �w  �uU  �8   �z�  ��  �h  Ӕ  ���|  �T  ���h  �T  ��$  ��  ���*  ��  ��y  �v  �  �u  �w  ��U   8   ���  X�  �h  Ӕ  ���|  �T  ���h  �T  ��$  X�  ���*  ]�  ��y  �v  �  �u  �w  �X  p�  ��  �h  l}  �j  �4&  ��   �b�  ev  @   ���  �  �p�  � �z�  ���  ���  @p5  ����  ���  � ���  @p5  ��ւ  ��̂  �    �SY  * �  6�  �h  ҡ  �4&  ��   ��  "�  `>   �R�  ��  ��  � �(�  ����  b�5  +��  �ւ  ��  �̂  �   ��T  ����Ge  �oY  / ��  ��  �h  ҡ  �-  �j  �4&  ��   ���  x~  �>   ���  _�  ���  � ���  ����  ����  ����  ��5  0D�  �ւ  A�  �̂  `�   ��T  ����Ge  ��Y  �   �w�  ��  �h  �  � �__s ���  ��ȱ  ���  ����� � ������  $u  ]u  ��Y  5�   ���  D�  �h  �  � �__s �D�  ��ȱ  �I�  ���j  ����� � ������  $u  ]u  ��Y   ,   �f�  ��  �h  �  ��__c �P(  ��w�  ��j  ��;�  ��j  ��__s ���  � 5y  �$Z  0   ���  �  �h  �  � �__c P(  ��;�� � ���  ��Z  @   � �  >�  �h  �  � ���  8>�  � 5y  �[  P   �[�  ��  �h  �  ��k  ����  T   C���  � �X�  T   	��}�  �p�  ��  �f�  �    m[   ��  ��  �h  �}  �__s P�j  |4&  P�   ���  �r  `�   ��  S�  ���  � ���  ��  ���  ��z6�  ��  ��3  ��ס  ��Ge  �[  a�  ��  �h  �~  �__s ��j  �4&  ��   �S�  d�  ��   ���  ��  �a�  � �k�  ��  �x�  ��
�L  �Z3  �p�xGe  �\  ��  �  �h  
�  �4&  c�   ���  �m  �>   �+�  ��  ���  � ��  ����  ��5  dg�  �ւ  ǧ  �̂  �   ��T  ����Ge  �\  ��  ��  �h  
�  �(�  q�-  �4&  q�   ���  �  �.   ���  "�  ���  � ���  �  ���  ����  �6  r�  �ւ  <�  �̂  [�   ��e   ��\  �   �:�  ��  �h  ��  � ���  ��j  ����  ��j  ����  ��j  ��k~  ��j  ����� � ������������  ��\   $   ���  �  �h  ��  ���k  ��j  ��:�  ��j  � �]  0   ��  j�  �h  ��  � ��k  ��j  ��:�  ��j  ��;�� � ������  �^  x�  ��  �h  ~  �__s  �j  �4&   �   �j�  n�  @�   ���  l�  �x�  � ���  z�  ���  ����  A06  9�  ��  ��  ���  ��  ���  A`6  d(�  �ւ  ��  �̂  ��   �dT  �� ��  ��3  ���  ��Ge ��Ge  v�c  ��e  �L   ���  �R  b  �ȱ  ���  � ��6  �__i ��c  N�  �E�  �{u  a�  ���  �'	�f �7	�i  �<	�f   ]u  L:  �  �  �h  �  �__c �q   ��R  @	�  �0�  ��  �h  ��  ��__s w�R  �  �$  w��  ���O  w�R  ��y  w�v  ���|  x�j  ��  ��h  x�j  � ��6  �ȱ  z��  ��w  {��  �  �}�  ]	   z��  ���  )�   ��6  ��  ��l  �q  �!�  �q  H�  �__c ��j  ��  ���  �	�6  �a�  ���  Ԫ  ���  �  ���  A�  ��6  �  u�    ���  �	7  ����  ��  ���  ��  ���  ݫ  �7  �  �  ���P   ���  �	87  }��  ���  �  ���  9�  ���  m�  �87  �  ��    ���  �
`7  ��  ��  ��  ��  ��  �n�  �
�7  ����  �  �|�  �  ��
!   x�  ���  P�z{  �
   ���{  ��{  !�    ��   ���  5�  �|�  �H��   ���  P    �n	r�    �u  ]u  l�  m7  ��  ��  �h  g�  }~�^  ��7  ~�&  �o6    J7  �  �  �h  g�  �__b ��   }y  �mW     �9�  ��  �h  Ӕ  ���|  J�T  ���h  J�T  �� �  J��  ���~  K�j  ���  K�j  � �R'  K�  �$�$  L��  �(��*  L��  �,��7  �ȱ  N��  ��w  O��  H�  �a�  R�j  g�  �__i U�  ��  �ȹ  V�j  ѭ  �}�  $   N<�  ���  �( ���  P�7  W��  ���  �  ��  F�7  ��,�  �  �F   ��  �7�  �{  O   B�+{  �5{  5�    � $   �,�  I�  � $   �7�      ���  `�7  W�  �ˆ  �$g  ���  �g  ���  `�7  ԍ�  �$g  ��  �g  �A�  `(8  �6�  �O�  �g  �(8  �Z�  ���  ``8  ��  ���  �g  �`8  ���  ���  \�  �F�  ��8  ��T�  Ϯ  ��    ��  �_�  ��  ��  �   V��  !�    �@	   �T�  4�  �@	   �_�  R�       ���  }�8  Ɲ��  p�  ���  (�     �A�  q�8  ��O�  �  ��8  �Z�  �  ���  q�8  Ɲ��  �  ��8  ���  �  ���  G�  �F�  w�8  ��T�  ��  �w   ��  �_�  ݱ  ��  �   V��  �    ��   �T�  *�  ��   �_�  >�           � 9  U�  �__c Y�j  ]�  �l�  �89  Y��  �z�  p�  ���  �89  ����  p�  �89  ���  ��  ���  ��  �F�  �`9  ��T�  \�  ��   ��  �_�  z�  ��  �   V��  ��    �h9  �T�  ��  �h9  �_�  Գ        ���  ��9  Y<�  ���  �  ���  �  ���  =�  ��9  �  ]�    ��9  �Р  ]�t  p�    ��  p   k��  ��  ��  ���  ��  ���  p   ���  ��  ���  ��    �1r�    �x  �u  �w  ]u  l�  �-W   X  ���  h�  �h  Ӕ  ���|  `�T  д  ��h  `�T  5�  �$  `h�  ���*  am�  ��y  a�v  � ��9  �ȱ  cr�  ��w  dw�  ���  e�j  �X��i  f�#  �\�}�  7   c��  ���  U�   �3�  ��9  o��  �[�  ��  �O�  ��  ���  ��9  Ν�  ��  ��  ��  �A�  ��9  ���  �O�  ��  ��9  �Z�  ۵  ���  �:  ���  ���  ��  �:  ���  ۵  ���  ��  �F�  �0:  ��T�  M�  ��   ��  �_�  k�  ��  �   V��  ��    �`	   �T�  V�`	   �_�  P     ���  �H:  Ɲ��  ��  ���  ��     �A�  �`:  ��O�  L�  �`:  �Z�  t�  ���  �`:  Ɲ��  L�  �`:  ���  t�  ���  ��  �F�   �:  ��T�  ݷ  �    ��  �_�  �   �	   �T�  �  �	   �_�  �           ��  �   p�  ��  �  ���  ,�  ���  �   ���  �  ���  @�    ��  �   mR�  ��  U�  ���  i�  ���  �   ���  U�  ���  }�    �@r�  �w!�    �u  �w  ]u  l�  v�e  ��e  �L   ���  �R  .\  �ȱ  ���  � ��:  �__i ��c  ��  �E�  �{u  ��  ���  ���f ���i  ���f   ]u  vi^  ��e  �L   ���  �R  D\  �ȱ  ���  � ��:  �__i ��c  ø  �E�  �{u  ָ  ���  ��f ��i  ��f   ]u  v�>  � f   L   ��  �R  1;  �ȱ  ��  � ��:  �__i ��c  ��  �E�  �{u  �  �-�  �W�f �g�i  �l�f   ]u  �>  pM  �)�  ��  �h  �  � �ȱ  N��  ���:  ��  ��#  R��  %�  ��  Tk  ��  ���  Uk  N�  ��  Vk  ,�  � ;  6�  ��b  o��  :�  �q�  �0;  Y��  ��  %�  �%�  �   ��3�  r�  ��  �Mz  �H;  YA�  �[z  ��  �4z  �   	��Bz  ��  �z  �   	-�$z  ��     ��  �`;  Y.�  ���  �  �4z  ��;  	#�  �Bz  �   ��}  ��;  	#��}  ��  ��}  #�  ��3   ��}  Y�  ��}  ��  �q}  ��;  	�!�  ��}  ��  �{}  ��  ��y  ��;  
V��y  ��  ��y  ��  ��;  �	z  Ǿ     ���     �q�  ��;  [o�  ��  ھ  �%�  �   ��3�  P�  �  ��  �;  [x�  ���  c�  �4z  <  	#��  �Bz  c�  �z     	-�$z  c�    ��}  &(<  	#��}  ӿ  ��}  C�  �P0   ��}  a�  ��}  ��  �q}  P@<  	�k�  ��}  ��  �{}  ��  ��y  P@<  
V��y  ��  ��y  ��  �@<  �	z  ��     �n�     ���  UX<  b��  ���  ��  �j�  e   ��x�  @�  �{  �Mz  ~   b�  �[z  S�  �4z  ~   	��Bz  S�  �z  ~   	-�$z  S�     ��  �p<  b��  ���  ��  �4z  �   	#N�  �Bz  ��   ��}  ��<  	#��}  M�  ��}  ��  �8��  �Rud   ���  ��<  d��  ���  ��  �j�  �   ��x�  S�  ��  ��  ��<  d?�  ���  q�  �4z  ��<  	#�  �Bz  q�   ��}  � =  	#��}  ��  ��}  ��  �H��  �Rud   ���  �=  g��  ���  ��  ���     ����  ��  �$  �Mz  '   g��  �[z  �  �4z  '   	��Bz  �  �z  '   	-�$z  �     ��  -0=  gN�  ���  ��  �4z  -   	#�  �Bz  ��   ��}  0P=  	#��}  D�  ��}  ��  ���  �Rud   ���  Sp=  i��  ���  ��  ���  c   ����  C�  �y  ��  ��=  i�  ���  V�  �4z  ��=  	#��  �Bz  V�   ��}  ��=  	#��}  ��  ��}  �  �(��  �Ru�   ���  ��=  lC�  �ϋ   �  ���  �   ���  >�    �ڋ  ��=  m~�  ��  Q�  �8�  �   ��F�  o�    ���  �>  p�  �Ʊ  ��  ���  ��  ���  ��  ���  �  �!�  5   ���  �S�  L�  �F�  _�  �9�  t�  �/�  ��   ���c   ���  J0>  s��  �Ʊ  ��  ���  ��  ���  ��  ���  ��  �!�  y+   �}�  �S�  1�  �F�  D�  �9�  Y�  �/�  l�   ���c   ��  �   [��  ���  ��  �4z  �   	#��  �Bz  ��   ��}  �   	#��}  ��  ��}  ��  ����  �Rud   ��  �!   ix�  ���  ��  �4z  �   	#=�  �Bz  ��   ��}  �   	#��}  ��  ��}  �  ����  �Ru�   ��  �   d��  ���  u\��4z  �   	#��  �Bz  u\� ��}  �   	#��}  �  ��}  K�  ����  �Rud   ��se �  ��se ��  �Gse ��  ��r�   ����  ���e ���e ���e ���d ��d �$�d �2�e �b�e �{�e  �kGe  ]u  ��  l�  v*M  �"f  �L   �7�  �R  G  �ȱ  �7�  � �X>  �__i ��c  ^�  �E�  �{u  q�  ���  ���f ��i  ��f   ]u  v G  �Df  L   ���  �R  U?  �ȱ  ���  � �p>  �__i ��c  ��  �E�  �{u  ��  ��  �G�f �W�i  �\�f   ]u  v3  �ff  `L   �E�  �R  �-  �ȱ  �E�  � ��>  �__i ��c  ��  �E�  �{u  ��  �m�  ���f ���i  ���f   ]u  ��2  ��  �b�  e �h  ��  � �ȱ  Ee ���>  Z �
m  Ij ��  ��  Pk  }�  �	v  Qk  ]�  ��p  Rk  ��  �ʌ  Sk  ��  ���  ��>  L�  ���  ��  �R�  �   ��`�  ��    ���  ��>  MN�  ���  ��  ���  �   ����  C�    �  �>  N��  �Њ  V�  �В     X�ޒ  ��    �?  � ��b  qo ��  �ۊ  H?  V��  ��  1�  ��  (   ��  ��  �>  �Mz  A   V;�  �[z  ��  �4z  A   	��Bz  ��  �z  A   	-�$z  ��     ��  G`?  V��  ���  g�  �4z  G   	#y�  �Bz  g�   ��}  J�?  	#��}  ��  ��}  ��  �x��  �Rud   �ۊ  m�?  X��  ��  ��  ��  }   ��  `�  ��  ��  ��?  Xj�  ���  ��  �4z  ��?  	#1�  �Bz  ��   ��}  ��?  	#��}  :�  ��}  ��  ����  �Rud   ��  �@  _��  ��  	�  �V�  �   &�d�  ��  �  �Mz     _�  �[z  ��  �4z     	��Bz  ��  �z     	-�$z  ��     ��  
 @  _y�  ���  o�  �4z  
   	#@�  �Bz  o�   ��}  @@  	#��}   �  ��}  ��  ���  �Rud   ��  0`@  a��  ��  ��  �V�  @   &�d�  {�  �V  ��  gx@  a1�  ���  ��  �4z  g�@  	#��  �Bz  ��   ��}  p�@  	#��}  !�  ��}  ��  �(��  �Rud   ��  ��@  dr�  ��  ��  ���  �   7���  '�  ��  �Mz  �   d��  �[z  P�  �4z  �   	��Bz  P�  �z  �   	-�$z  P�     ��  ��@  d@  ���  ��  �4z  �   	#  �Bz  ��   ��}  � A  	#��}  ��  ��}  <�  �X��  �Rud   ��  � A  f�  ��  Z�  ���  �   7���  ��  ��  ��  8A  f�  ���  �  �4z  XA  	#�  �Bz  �   ��}  pA  	#��}  ��  ��}  2�  �h��  �Rud   �&�  '�A  i9 �4�  P�  ���  7   H��  ��  �P  �Mz  S   i� �[z  ��  �4z  S   	��Bz  ��  �z  S   	-�$z  ��     ��  Y�A  i ���  1�  �4z  Y   	#� �Bz  1�   ��}  \�A  	#��}  ��  ��}  ��  �8��  �Rud   �&�  �A  kH �4�  �  ���  �   H��  I�  ��  ��  ��A  k� ���  \�  �4z  �B  	#� �Bz  \�   ��}  �0B  	#��}  ��  ��}  �  �H��  �Ru�   �?�  �HB  n� �M�  &�  ��  �   |��  D�    �X�  �`B  o7 �f�  W�  �N�  �   ��\�  u�    ���  xB  r� �Ʊ  ��  ���  ��  ���  ��  ���  ��  �!�  7   �� �S�  "�  �F�  5�  �9�  J�  �/�  ]�   �k�c   ��     a3 ���  �  �4z     	#� �Bz  �   ��}     	#��}  ��  ��}  ��  �!��  �Rud   ��  ^   X� ���  ��  �4z  ^   	#q �Bz  ��   ��}  d   	#��}  ��  ��}  �  �s��  �Rud   ��  �)   k# ���  )�  �4z  �   	#� �Bz  )�   ��}  �#   	#��}  >�  ��}  S�  ����  �Ru�   ��  �B   f� ���  f�  �4z  �   	#a �Bz  f�   ��}  �<   	#��}  {�  ��}  ��  �
 ��  �Rud   �ase ��  �$se �g  ��se �  �sse ��  �r�   ����  ���e ���d ���d ���d ��d ��e �M�e �|�e ���e  �VGe  ]u  ��  l�  v�-  ��f  @ L   �� �R  �(  �ȱ  �� � ��B  �__i ��c  ��  �E�  �{u  ��  �M �  �w �f �� �i  �� �f   ]u  �d-  � �  �  �h  �  � �ȱ  E ���B   �
m  I ��  ��  Pk  x�  �	v  Qk  X�  ��p  Rk  ��  �ʌ  Sk  ��  ���  � �B  L� ���  ��  ��  �    ��%�  ��    ���  � �B  M� ���  ��  �V�  �    ��d�  >�    ���  � C  N: �ǉ  Q�  ���  �    X���  ��    � C  � ��b  q  ��  �҉  � `C  V� ���  ,�  ���  !   ��  ��  �!  �Mz  !!   V� �[z  ��  �4z  !!   	��Bz  ��  �z  !!   	-�$z  ��     ��  '!xC  Vc	 ���  b�  �4z  '!   	#*	 �Bz  b�   ��}  *!�C  	#��}  ��  ��}  ��  �X&��  �Rud   �҉  M!�C  X�	 ���  ��  ���  ]!   ��  [�  �s!  ��  �!�C  X
 ���  ��  �4z  �!�C  	#�	 �Bz  ��   ��}  �!D  	#��}  5�  ��}  ��  �h&��  �Rud   ��  �! D  _\
 ��  �  �B�  �!   &�P�  ��  ��!  �Mz  �!   _�
 �[z  ��  �4z  �!   	��Bz  ��  �z  �!   	-�$z  ��     ��  �!8D  _* ���  j�  �4z  �!   	#�
 �Bz  j�   ��}  �!XD  	#��}  �  ��}  ��  ��%��  �Rud   ��  "xD  ak ��  ��  �B�   "   &�P�  v�  �6"  ��  G"�D  a� ���  ��  �4z  G"�D  	#� �Bz  ��   ��}  P"�D  	#��}  �  ��}  ��  �&��  �Rud   �'�  a"�D  d# �5�  ��  ���  q"   7���  "�  ��"  �Mz  �"   dz �[z  K�  �4z  �"   	��Bz  K�  �z  �"   	-�$z  K�     ��  �"�D  d� ���  ��  �4z  �"   	#� �Bz  ��   ��}  �"E  	#��}  ��  ��}  7�  �8&��  �Rud   �'�  �"8E  f2 �5�  U�  ���  �"   7���  ��  ��"  ��  �"PE  f� ���  ��  �4z  �"pE  	#p �Bz  ��   ��}  �"�E  	#��}  ��  ��}  -�  �H&��  �Rud   �@�  #�E  i� �N�  K�  �̘  #   H�ژ  ��  �0#  �Mz  3#   iA �[z  ��  �4z  3#   	��Bz  ��  �z  3#   	-�$z  ��     ��  9#�E  i� ���  ,�  �4z  9#   	# �Bz  ,�   ��}  <#�E  	#��}  ��  ��}  ��  �&��  �Rud   �@�  _#�E  k� �N�  �  �̘  o#   H�ژ  D�  ��#  ��  �#F  kr ���  W�  �4z  �#0F  	#7 �Bz  W�   ��}  �#HF  	#��}  ��  ��}  �  �(&��  �Ru�   �Y�  �#`F  n� �g�  !�  �ԑ  �#   |��  ?�    �r�  �#xF  o� ���  R�  ��  �#   ��!�  p�    ���  �#�F  rm �Ʊ  ��  ���  ��  ���  ��  ���  ��  �!�  $   �b �S�  �  �F�  0�  �9�  E�  �/�  X�   �K$�c   ��  �&   a� ���  z�  �4z  �&   	#� �Bz  z�   ��}  �&   	#��}  ��  ��}  ��  �'��  �Rud   ��  >'   X[ ���  ��  �4z  >'   	#" �Bz  ��   ��}  D'   	#��}  ��  ��}  �  �S'��  �Rud   ��  �')   k� ���  $�  �4z  �'   	#� �Bz  $�   ��}  �'#   	#��}  9�  ��}  N�  ��'��  �Ru�   ��  �'B   fK ���  a�  �4z  �'   	# �Bz  a�   ��}  �'<   	#��}  v�  ��}  ��  ��'��  �Rud   �A!se ��!  �"se �G"  ��"se ��"  �S#se ��#  ��#r�   �� z ��&�e ��&�d ��&�d ��&�d ��&�d ��&�e �-'�e �\'�e ��'�e  �6'Ge  ]u  t l�  v,;  ��f   (L   �� �R  �7  �ȱ  �� � ��F  �__i ��c  ��  �E�  �{u  ��  �-(�  �W(�f �g(�i  �l(�f   ]u  v�7  ��f  p(L   �. �R  4  �ȱ  �. � ��F  �__i ��c  ��  �E�  �{u  ��  �}(�  ��(�f ��(�i  ��(�f   ]u  v�R  ��f  �(L   �� �R  :M  �ȱ  �� � ��F  �__i ��c    �E�  �{u  +  ��(�  ��(�f �)�i  �)�f   ]u  �:  � � �h  �  ��+  �j  �R'  /M   ��S  )�  �  �h  ��  ��__s ��R  I  �$  � ���R  ��y  ��v  ���l  �q  ��!�  �q  � � G  �ȱ  � ��w  � }  �'y  � �  �ǆ  ��c  ��/t  �# ��~�-  �Zw  ��~�}�  4)   �� ���  �   ��  T)G  �< ���  %��  �  �`*E   ���  %��  V�o*�c    ��  �)8G  �\ ���    ��  �)XG  �� �5�  > �*�  Q ��  u �� �)pG  r�� > �� Q �� � ���  �)   ��  � �؅   �΅  "    �F)r�  �T)9 ��)�M    �u  ]u  l�  3 wq  3 z)l   v�S  �g  �*L   �� �R  �R  �ȱ  �� � ��G  �__i ��c  5 �E�  �{u  H ��*�  ��*�f ��*�i  ��*�f   ]u  v�X  �2g   +L   �< �R  MT  �ȱ  �< � ��G  �__i ��c  f �E�  �{u  y �+�  �7+�f �G+�i  �L+�f   ]u  vK[  �Tg  P+L   �� �R  �X  �ȱ  �� � ��G  �__i ��c  � �E�  �{u  � �]+�  ��+�f ��+�i  ��+�f   ]u  �vg  �+I   �4 �R  b  �ȱ  h4 � ��+@   �__i j�c  � �E�  k{u  � ��+�  ��+�f   ]u  ��g  �+I   �� �R  .\  �ȱ  h� � ��+@   �__i j�c  � �E�  k{u   ��+�  �,,�f   ]u  ��g  @,I   � �R  D\  �ȱ  h � �D,@   �__i j�c  * �E�  k{u  H �N,�  �|,�f   ]u  ��g  �,I   �� �R  1;  �ȱ  h� � ��,@   �__i j�c  [ �E�  k{u  y ��,�  ��,�f   ]u  ��g  �,I   �� �R  G  �ȱ  h� � ��,@   �__i j�c  � �E�  k{u  � ��,�  �-�f   ]u  � h  0-I   �i �R  U?  �ȱ  hi � �4-@   �__i j�c  � �E�  k{u  � �>-�  �l-�f   ]u  �Bh  �-I   �� �R  �(  �ȱ  h� � ��-@   �__i j�c  � �E�  k{u   ��-�  ��-�f   ]u  �dh  �-I   �K �R  �7  �ȱ  hK � ��-@   �__i j�c   �E�  k{u  = ��-�  �.�f   ]u  ��h   .I   �� �R  4  �ȱ  h� � �$.@   �__i j�c  P �E�  k{u  n �..�  �\.�f   ]u  ��h  p.I   �- �R  :M  �ȱ  h- � �t.@   �__i j�c  � �E�  k{u  � �~.�  ��.�f   ]u  ��h  �.I   �� �R  �R  �ȱ  h� � ��.@   �__i j�c  � �E�  k{u  � ��.�  ��.�f   ]u  ��h  /I   � �R  MT  �ȱ  h � �/@   �__i j�c  � �E�  k{u   �/�  �L/�f   ]u  �i  `/I   �� �R  �X  �ȱ  h� � �d/@   �__i j�c   �E�  k{u  2 �n/�  ��/�f   ]u  �0i  �/�  �g !T  q  �__s �k  E �3�  �q  ���  ��j  ��V�  ��  ��z  ��j   ��l  ��j  � ��G  ��p  ��  � ���  ��  E ��G  I �__i �q  �  ��0<   �__i �q  �    ��H  `1�   � �  �h  ]�  � ��  ��j  ����  ��  ��3�  �q  ��__p ��j  ���  �k  ����  �k  ��R'  ��  ��H  ���  ��t  � �ʞ  �k  ' ��l  ��j  E ��  �1 H  �s  ��  n ��  � ��  � ��1#e  ��1� ��1�   �x  �5I   25   ��  C! �h  ]�  � ��  B�j  ����  B�  ��3�  Bq  ��C! ���  Ck  ����  Ck  ��R'  CH! ��2   �__p Ek  � �+2�   �u  �x  �`  [! �! �h  �! |ȱ  +�! }�__i -�c  ~C�  .{u  }~Y�  1�w     �y  ]u  j  �! �! �h  %~  �%  	d�  �__n 	d�     �! " �h  %~  �%  	9�  �__n 	9�  �__c 	9q   �A9  @2  �6" �. Y�  �t  �h  �  ��__s ��7  � �$  ��. ���O  ��7  ��{�  ��. ��8H  q. T�e  ��  T�k  ��'  T��  ��1  �ȱ  ��. ��w  ��. � �ϴ  ��`  ��k  ��" �" �" �ԥ  ��. ��|  ��. J	 �__p ��'  �\�gh  ��. �	 �x  ��" �	 �R'  ��" 
 �}�  e2PH  �v# ���  �
  �M! t2hH  �r$ �e! �
 �[! �  �hH  �q! - �}! l ��H  f$ ��! � ���  �8|   4$ ���  � ���   ���  �8   ��ւ  � �̂     ��8g �s9J�  ��9�  �3:�e �;:�e �D:�e �U:�e  ��2�    �T�  �2   ��$ �b�  : �z  �2   	&�$z  :   �}�  �2�H  ��% ���  f ���  � ���  	 ���  M ��H  ���  ���  y ���  ���  ��   6�H  ��3�  � �'�   ��  ��H  ��  �3�  � �'�   ��H  �@�  2 �K�  �V�  � �I  �b�  Z �HI  �n�  � ��6f ��7�e �>8�f �^8�e �~8af ��8Lf ��87f        �xI  . �ȹ  �8  �T��p  �%   ` �__f ��$  �/t  �8  �X�8w  �=& � �" �S�  �u   ���  $3   ��& ���  N �X�  $3   	��}�  �p�  � �f�     ��I  ) ��  �k  � �m�  b3�I  �' ���  � ���   �{�  � �Mz  j3   	�' �[z  �  �{3h   ��  �3�I  ��' ��  � ���  � �~  �3�I  	\�~  � �4z  �3   	<�' �Bz  � �z  �3   	-�$z  �   ��3�	    ��  �3�I  �0( ��  3 ���  S �~  �3�I  	\�~  S �4z  �3   	<$( �Bz  S �z  �3   	-�$z  S   ��3�	    ��! �3J  �) ��! � ��! � ��! � �*~  �3   	g�( �O~  � �B~  � �8~  � ��3   �]~   �Mz  �3   	U�[z  �    �l~  �3 J  	g) ��~  ' ��~  O �z~  m ��9�i   �4�	   ��3�  ���  48J  �P) �Ȍ  � ���  � �(4��   �(�  K4PJ  �z) �>�  3 �2�  |  ���  {4   ��) ���  � �X�  {4   	��}�  �p�  � �f�  �   �xJ  �* �__i ��j   ��J  ���  ��) � �" ���  7   1* �Ȍ  ) ���  > �7��   ���  @7   e* ���  S ���  � �M7�   ���  �9   �* �Ȍ  ���  � ��9��   ��6�  �77&    �Mz  
5   + �[z  � �4z  
5   	��Bz  � �z  
5   	-�$z  �    ��! #5�J  #K+ �" � ��! � ��!  ��! 3 �;5h   ��  A5�J  (�+ �5�  H �*�  s ��  � �� A5�J  r�� H �� s �� � ���  G5   ��   �؅  ! �΅  4    ��  f5�J  �V, ���  T �4z  f5   	#, �Bz  T  ��}  i5K  	#��}  v ��}  � ��9��  �Ru[   ��  t5   (�, ���  � �4z  t5   	#�, �Bz  �  ��}  z5   	#��}  � ��}  � ��5��  �Rw    ��  �9   �F- ���  � �4z  �9   	#- �Bz  �  ��}  �9   	#��}   ��}  5 �:��  �Ru[   ��  :   (�- ���  H �4z  :   	#�- �Bz  H  ��}  :   	#��}  ] ��}  � �!:��  �Ru`   �533  �H4�  ��43  �5�  �p7�  ��7&  ��7�  ��9&   ���  �5(K  *F. ���  ���  � �(K  �ρ  �   �Mz  �5   �f. �[z  �  �t2r�   �*:Ge �^:Ge  �u  x  ]u  l�  ~9  8a  �. �. �h  �. |ȱ  +�. }�__i -�c  ~C�  .{u  }~Y�  1�w     �y  ]u  ��9  `:  �/ f; Y�  �t   �h  �  ��__s ��7  � �$  �f; ���O  ��7  ��{�  �k; ��@K  Q; T�e  ��  T�k  ��'  T��  �B,  �ȱ  �p; ��w  �u;  �ϴ  �,a  ��k  ��/ �/ �/ �ԥ  ��. ��|  ��. P �__p ��'  �\�gh  ��. � �x  �n/ � �R'  �n/  �}�  �:XK  �V0 ���  �  ��. �:pK  �R1 ��. � ��. �~�  �pK  ��. 3 ��. r ��K  F1 ��. � ��  A|   4�0 �7�  � �-�   ���  A   ��ւ  � �̂     �
Ag ��A� ��A�  �SB�e �[B�e �dB�e �uB�e  ��:�    �T�  �:   ��1 �b�  @ �z  �:   	&�$z  @   �}�  �:�K  ��2 ���  l ���  � ���    ���  S  ��K  ���  ���    ���  ���  ��  @>�K  ��3�  �  �'�  ! ��  ��K  ��  �3�  �  �'�  ! ��K  �@�  8! �K�  �V�  �! � L  �b�  `" �PL  �n�  �" ��>f �@�e �^@�f �~@�e ��@af ��@Lf ��@7f        ��L  �: �ȹ  �8  �T��p  �%   f# �__f ��$  �/t  �8  �X�8w  �3 �# n/ �S�  �u  $ ���  D;   �3 ���  T$ �X�  D;   	��}�  �p�  �$ �f�  %   ��L  �5 ��  �k  �% �m�  �;�L  ��3 ���  �% ���  & �{�  �& �Mz  �;   	��3 �[z  �&  ��;h   ��  �;�L  ��4 ��  �& ���  �& �~  �;�L  	\�~  �& �4z  �;   	<x4 �Bz  �& �z  �;   	-�$z  �&   ��;�	    ��  �;�L  �5 ��  9' ���  Y' �~  �;�L  	\�~  Y' �4z  �;   	<5 �Bz  Y' �z  �;   	-�$z  Y'   �<�	    ��! <M  ��5 ��! �' ��! �' ��! �' �*~  <   	g�5 �O~  �' �B~  �' �8~  �' �<   �]~  ( �Mz  <   	U�[z  �'    �l~  <(M  	g�5 ��~  -( ��~  U( �z~  s( �B�i   �'<�	   ��;�  ���  4<@M  �06 �Ȍ  �( ���  �( �H<��   �(�  k<XM  �Z6 �>�  9) �2�  �)  ���  �<   ��6 ���  �) �X�  �<   	��}�  �p�  �) �f�  �)   ��M  �7 �__i ��j  * ��M  ���  ��6 �* z/ ���  &?   7 �Ȍ  /+ ���  D+ �2?��   ���  `?   E7 ���  Y+ ���  �+ �m?�   ���  �A   u7 �Ȍ  ���  �+ ��A��   �?�  �W?&    �Mz  *=   �7 �[z  �+ �4z  *=   	��Bz  �+ �z  *=   	-�$z  �+    ��! C=�M  #+8 �" �+ ��! , ��! %, ��! 9, �[=h   ��  a=�M  (�8 �5�  N, �*�  y, ��  �, �� a=�M  r�� N, �� y, �� �, ���  g=   ��  - �؅  '- �΅  :-    ��  �= N  �69 ���  Z- �4z  �=   	#�8 �Bz  Z-  ��}  �=N  	#��}  |- ��}  �- ��A��  �Ru[   ��  �=   (�9 ���  �- �4z  �=   	#u9 �Bz  �-  ��}  �=   	#��}  �- ��}  �- ��=��  �Rw    ��  B   �&: ���  �- �4z  B   	#�9 �Bz  �-  ��}  B   	#��}  . ��}  ;. �,B��  �Ru[   ��  ,B   (�: ���  N. �4z  ,B   	#e: �Bz  N.  ��}  2B   	#��}  c. ��}  �. �AB��  �Ru`   �U;3  �h<�  ��<3  �'=�  ��?�  ��?&  ��?�  ��A&   ���  �=0N  *&; ���  ���  �. �0N  �ρ  �.   �Mz  �=   �F; �[z  �.  ��:r�   �JBGe �~BGe  �u  x  ]u  l�  ��8  �B�  ��; p? �h  �  ��__s :�7  ����  :�t  ��$  :p? ���O  :�7  ��#�  ;st  ��HN  e? �ȱ  =�!  �X��w  >u? �. ���  Q�t  / ���  Sk  :/ �R'  T�j  r/ �{�  W8  �\�ˍ  �BhN  =�< �ٍ  ���B ��  �B�N  X= ��  �/ ���  �/ �~  �B�N  	\�~  �/ �4z  �B�N  	<= �Bz  �/ �z  �B�N  	-�$z  �/   �C�	    ���  C�N  X�= �Ʊ  0 ���  .0 ���  I0 ���  ^0 �!�  :C   ��= �S�  |0 �F�  �0 �9�  �0 �/�  �0 �KC#e  ��C�c   ��  qC�N  W�> ���  �0 �4z  qC�N  	#�= �Bz  �0 �z  qC   	-�$z  �0   ��}  zCO  	#��}  1 ��}  E1 � D.   ��}  c1 ��}  �1 �q}   D(O  	��> ��}  �1 �{}  �1 ��y   D(O  
V��y  �1 ��y  �1 �(O  �	z  �1    �D�     ��  .D   W ? ���  �1 �4z  .D   	#�> �Bz  �1  ��}  4D   	#��}  2 ��}  /2 �CD��  �R�W   ��Br�  ��BT  ��B��  ��B�qC" ��C��C�. �LD �TDGe  �u  l�  �9  `Dw   ��? @ �h  �  ��__s `�7  ����  `�t  ��$  `@ ���O  `�7  ��{�  a	@ ���D�. ��D"  �u  x  ��^  �D4  �C �$  �C � ��O  �q  ����  �k  B2 �A�  ��j  ���l  �/M  ��G�  �/M  ��@O  ���  ��c  �2 ��h  ��$  �!�  ��   3 �(�  EhO  ��@ �>�  ��2�  g3  ��O  �B �ȱ  ��C ��w  ��C �3 �}�  cE   �'A ���  �3  ��  lE�O  �vA ���  4 ��  �3 ��O  ���  ;4 ��  ]4 �-F�c    ��  �E�O  ��A ���  �4 ��  �4 ��F_�  �P�\�RX  ��  UF   ��A ���  �4 ��  �4 �oF_�  �P�\�R+  ��  �F   �BB ���  "5 ��  Q5 ��F_�  �P�\�R0  ��  �F   ��B ���  {5 ��  �5 ��F_�  �P�\�Rx  �lEr�   �K�  !E�O  ��B �o�  �5 �b�  �5 �U�  6 �3E g  ��  7EP  �	C ��  !6 ��  c6 ��  �SE#e  ��  �E0P  �GC ��  �6 ��  �6 ��  �6 ��E#e  �K�  �EHP  ��o�  7 �b�  7 �U�  ��E g    �u  ]u  l�  �sI   G/   ��C D �h  ]�  � ��O  q  ��__w /M  ��$  D ���  k  ����  �j  ��R'  #D ��GG@  �u  �x  �li  PG�   �+E !T  q  ]T  7   �{�  k  G7 �__v 7   }7 �ԥ  �j  �7 ���  �#  ����  �t  ��`P  ���  k  8 �(�  �G   #�D �>�  J�2�  � ��P  ���  0u  _8 ��j  1�t  �(�  �G�P  0�>�  �8 �2�  �8     ua  9E uE �h  uE |ȱ  5zE }�__i 7�c  ~C�  8{u  }~Y�  ;Sx     �y  ]u  ��K   H  ��E qI ]T  %   �h  ]�  ��__s N�9  �8 �$  NqI ���O  Nq  ��__v O%   ���P  fI Tߠ  R�l  T��  S�=  �ϴ  Tia  �ȱ  UvI ��k  V7F =F F �ԥ  W�j  �8 ���  X�$  ���  [�t  9 ���  \k  19 ��m  a�$  ���  bu  d: �__u d�F �: �E �R'  g�j  �\�__w ��i  �+E H�P  V�G �CE ; �9E ���  ��P  �OE N; �[E �; �Q  �G �gE �; ��  QJ0Q  >|G ��  �; ��   < ���  QJ   ?�ւ  �; �̂   <   �JJg ��J�  ��J�  ��J�e ��J�e ��J�e ��J�e  �%H�    �(�  VHHQ  a�G �>�  I< �2�  k<  ��ID   #H ���  ok  �< ��I�   ��I6   CH ���  �u  �<  ��H/   mH ���  �k  �< �I�C  ���  I   ��H ���  ���  �< �I   �ρ  �<   ��  I2   �;I �5�  = �*�  "= ��  5= �� I#   r�� = �� "= �� �= ���  $I   ��  �= �؅  �= �΅  �=    �}�  MJhQ  U[I ���  �=  ��H(D  �KGe  �u  ]u  ��I  K�  ��I �O �h  ]�  ��__s A6G  $> �$  A�O ���O  A)G  ��__v A�t  ���Q  �O ���  C�$  �(�  /K�Q  DJ �>�  �2�  8>  ��Q  EJ �__l F�y  o> �ZKE  ��Q  T��  K�=  �ϴ  Lia  �ȱ  M�O ��k  N~J �J KJ �F�  P�j  �> �R'  R�j  �> �__w U�i  �+E �K R  N�K �CE "? �9E �%�  � R  �OE t? �[E �? �(R  �K �gE �? ��  DMG   >aK ��  P@ ��  |@ ���  DM   ?�ւ  P@ �̂  |@   �:Mg ��M�  ��M�  ��M�e ��M�e ��M�e ��M�e  ��K�    �HR  �N ���  X�i  �@ ��  Yk  �@ �K�  �KpR  ]L �o�  �A �b�  �A �U�  �@ ��K g  �(�  �K�R  `HL �>�  �A �2�  .B  ���  L   ^�L ���  ZB ���  �B �L   �ρ  �B   ��   L�R  gM �5�  �B �*�  �B ��  �B ��  L�R  r�� �B �� �B �� C ���  )L   ��  +C �؅  >C �΅  QC    ��  BL   h�M �5�  dC �*�  �C ��  �� BL   r�� dC �� �C �� �C ���  BL   ��  dC �؅  �C �΅  �C    ��  �L+   b<N �5�  �C �*�  �C ��  D �� �L+   r�� �C �� �C �� +D ���  �L   ��  CD �؅  nD �΅  �D    ��  M%   c�5�  �D �*�  �D ��  �� M%   r�� �D �� �D �� �D ���  M   ��  �D �؅  �D �΅  �D     ��  �L�R  m[O �5�  �D �*�  E ��  %E �� �L�R  r�� �D �� E �� OE ���  �L   ��  gE �؅  �E �΅  �E    ���  �L   l�O ���  �E ���  �E ��L   �ρ  �E   �}�  =M   M���  �E    ��MGe  �u  ]u  J  �O P �h  ]�  �__s �	6G  �$  �	P ��O  �	)G  �__v �	%    �u  ��O �s   N1   �;P sP ��O ���O ���O ���O ��P ��(NE  ��G  @Nr   ��P #Q �h  ]�  ��__s 	6G  ��$  	#Q ���O  	)G  ��__v 	%   ���O cN    	�P )F ��O =F ��O QF ��O ��O pF �{NE   �u  ��K  �N�  �IQ U ]T  7   �h  ]�  ��__s N�9  �F �$  NU ���O  Nq  ��__v O7   ���R  U Tߠ  R�s  T��  S�=  �ϴ  Tia  �ȱ  UU ��k  V�Q �Q �Q �ԥ  W�j  �F ���  X�$  ���  [�t  G ���  \k  ,G ��m  a�$  ���  bu  �G �__u dZR �G �Q �R'  g�j  �\�__w ��i  �+E �N�R  VxS �CE �G �9E ��  ��R  �OE EH �[E yH �(S  lS �gE �H ��  �PG   >%S ��  �H ��  "I ���  �P   ?�ւ  �H �̂  "I   ��Pg ��P�  �Q�  �-Q�e �=Q�e �FQ�e �OQ�e  ��N�    �(�  OHS  a�S �>�  VI �2�  xI  �`S  �S ���  ok  �I �+P�   �aP/   �S ���  �u  �I  �wO1   T ���  �k  �I ��O�C  ���  �O   �MT ���  ���  �I ��O   �ρ  J   ��  �O,   ��T �5�  *J �*�  =J ��  PJ �� �O!   r�� *J �� =J �� �J ���  �O   ��  �J �؅  �J �΅  �J    �}�  �P   U U ���  K  �IO(D  �XQGe  �u  ]u  CJ  .U mU �h  ]�  �__s �	6G  �$  �	mU ��O  �	)G  �__v �	7    �u  � U ��  `Q1   ��U �U �.U ��8U ��EU ��RU ��_U ���Q(Q  �jK  �Qp   ��U �V �h  ]�  ��__s �6G  ?K �$  ��V ���O  �)G  ��__v �l  ���QL   ���  ��$  �-  ��$  �(�  �Q   �yV �>�  ��~�2�  cK  ��  �Q   ��V �4�  �(�  �K  �=�  �Q   ��V �K�  �K �U�  �K ��Q   �c�    ��Q(Q   �u  ��G  Rr   �W �W �h  ]�  ��__s #	6G  ��$  #	�W ���O  #	)G  ��__v $	7   �� U 3R   %	�_U L �RU $L �EU 8L �8U �.U WL �KR(Q   �u  ��i  �R  ��X !T  q  ]T  )k  �{�  k  � �__v )k  vL �ԥ  �j  ����  �#  ����  �t  ��xS  ���  k  �L �(�  
S   #VX �>�  J�2�  � ��S  ���  0u  CM ��j  1�t  �(�  S�S  0�>�  �M �2�  �M     �L  �S(  ��X �\ ]T  0k  �h  ]�  ��__s N�9  �M �$  N�\ ���O  Nq  ��__v O0k  ���S  �\ Tߠ  R�l  T��  S�=  �ϴ  Tia  �ȱ  U�\ ��k  V[Y aY (Y �ԥ  W�j  �M ���  X�$  ���  [�t  N ���  \k  @N ��m  a�$  ���  bu  sO �__u d�Y �O Y �R'  g�j  �\�__w ��i  �+E �S�S  V�Z �CE �O �9E ��  ��S  �OE �O �[E P �(T  �Z �gE @P ��  !VPT  >�Z ��  �P ��  �P ���  !V   ?�ւ  �P �̂  �P   �Vg �rV�  ��V�  ��V�e ��V�e ��V�e ��V�e  ��S�    �(�  ThT  a[ �>�  �P �2�  Q  ��T  C[ ���  ok  @Q �U�   ��U8   c[ ���  �u  `Q  ��T2   �[ ���  �k  }Q ��T�C  ���  �T   ��[ ���  ���  �Q ��T   �ρ  �Q   ��  �T*   �[\ �5�  �Q �*�  �Q ��  �Q �� �T   r�� �Q �� �Q �� #R ���  �T   ��  ;R �؅  NR �΅  aR    �}�  V�T  U{\ ���  uR  �pT�W  ��VGe  �u  ]u  ~J  �\ �\ �h  ]�  �__s �	6G  �$  �	�\ ��O  �	)G  �__v �	0k   �u  ��\ >�  �V5   �	] A] ��\ ���\ ���\ ���\ ���\ ��W�X  ��G   Wo   �Y] �] �h  ]�  ��__s )	6G  ��$  )	�] ���O  )	)G  ��__v )	0k  ���\ MW   *	��\ �R ��\ �R ��\ �R ��\ ��\ �R �`W�X   �u  �YL  �W�  �^ �a ]T  )k  �h  ]�  ��__s N�9  S �$  N�a ���O  Nq  ��__v O)k  ���T  �a Tߠ  R�s  T��  S�=  �ϴ  Tia  �ȱ  U�a ��k  V�^ �^ {^ �ԥ  W�j  \S ���  X�$  ���  [�t  �S ���  \k  �S ��m  a�$  ���  bu  2T �__u d(_ qT o^ �R'  g�j  �\�__w ��i  �+E �W�T  VF` �CE �T �9E �U�  ��T  �OE �T �[E U �U  :` �gE 2U ��  �Y0U  >�_ ��  U ��  �U ���  �Y   ?�ւ  U �̂  �U   ��Yg ��Y�  ��Y�  �Z�e �-Z�e �6Z�e �?Z�e  ��W�    �(�  �WHU  ap` �>�  �U �2�  �U  ��XF   �` ���  ok  0V �Y�   �GY9   �` ���  �u  aV  �VX1   �` ���  �k  }V �X�C  ���  �X   �a ���  ���  �V ��X   �ρ  �V   ��  �X,   ��a �5�  �V �*�  �V ��  �V �� �X!   r�� �V �� �V �� FW ���  �X   ��  ^W �؅  qW �΅  �W    �}�  �Y`U  U�a ���  �W  �(X�W  �HZGe  �u  ]u  �J   b ?b �h  ]�  �__s �	6G  �$  �	?b ��O  �	)G  �__v �	)k   �u  ��a �f  PZ5   �`b �b � b ��
b ��b ��$b ��1b ��|Z�]  �+H  �Zo   ��b Hc �h  ]�  ��__s -	6G  ��$  -	Hc ���O  -	)G  ��__v .	)k  ���a �Z   /	�1b �W �$b �W �b �W �
b � b X ��Z�]   �u  �M! W�   [(  �ic Yd �[! � �e! ��xU  Nd �q! :X �}! nX ��U  Cd ��! �X ���  L[|   4�c ���  Y ���  GY ���  L[   ��ւ  Y �̂  GY   �J[g ��[J�  ��[�  ��[�e �\�e �\�e �\�e  �[�   �(\Ge  ��. ��  0\(  �ud ee ��. � ��. ���U  Ze ��. �Y ��. �Y ��U  Oe ��. Z ��  |\|   4e �7�  kZ �-�  �Z ���  |\   ��ւ  kZ �̂  �Z   �z\g �]� �]�  �*]�e �2]�e �;]�e �O]�e  �F\�   �X]Ge  �+E ��  `]�   ��e qf �9E � �CE ���U  ff �OE �Z �[E [ �V  [f �gE T[ ��  �]G   >f ��  �[ ��  �[ ���  �]   ?�ւ  �[ �̂  �[   ��]g ��]�  �^�  �%^�e �-^�e �6^�e �J^�e  �v]�   �S^Ge  ��L  `^�  ��f \j ]T  zt  �h  ]�  ��__s ��9  *\ �$  �\j ���O  �q  ��!�  �q  ��__v �zt  �� V  T��  ��=  �ϴ  �ia  �G�ȱ  �aj ��k  �0g o\ 6g �f ��6  ��i  �\ �+w  ��t  �R'  ��j  �H�w  �fj �P��  �u  �\ �4�  ��t  4���  ��t  �\ ���  �k  ] ��w  vj ;] ��+  k  q] ��  
k  �] �__p �j  �__w /�i  �}�  �^   �)h ���  �]  ���  +_PV  �h �Ʊ  ^ ���  .^ ���  f^ ���  �^ �!�  Q_   ��h �S�  �^ �F�  �^ �9�  �^ �/�  �^_#e  ��`�c  �0a#e  �I  f_   �h �m  �`  _ �S  V_ �u_Bg  �xV  0i ��  k  _ �Q  /M  �_ ��`g  ��_5   Zi �0�  2k  �_ ��_�C  ���  �_   7�i ���  ���  �_ ��_   �ρ  �_   ��  �_4   ;(j �5�  ` �*�  2` ��  G` �� �_)   r�� ` �� 2` �� �` ���  �_   ��  �` �؅  �` �΅  �`    ��^+E ��^�&  ��^T  �_��  �_r�    �u  ]u  wq  vj z)l   l�  ��J  @a7   ��j �j �h  ]�  ��__s u6G  ��$  u�j ���O  u)G  ��__v uzt  ��naqf  �u  ��L  �a�  �k �n ]T  st  �h  ]�  ��__s ��9  a �$  ��n ���O  �q  ��!�  �q  ��__v �st  ���V  T��  ��=  �ϴ  �ia  �G�ȱ  ��n ��k  ��k Xa �k uk ��6  ��i  �a �+w  ��t  �R'  ��j  �H�w  �fj �P��  �u  �a �4�  ��t  D���  ��t  �a ���  �k  �a ��w  �n $b ��+  k  Zb ��  
k  �b �__p �j  �__w /�i  �}�  �a   ��l ���  �b  ���  Eb�V  >m �Ʊ  �b ���  ec ���  �c ���  �c �!�  kb   �)m �S�  d �F�  d �9�  4d �/�  �xb#e  ��c�c  �Pd#e  �I  �b   xm �m  �`  Gd �S  �d ��bBg  ��V  �m ��  k  �d �Q  /M  �d ��cg  ��b5   �m �0�  2k  e ��b�C  ���  �b   7n ���  ���  !e ��b   �ρ  5e   ��  �b4   ;�n �5�  Ie �*�  ie ��  ~e �� �b)   r�� Ie �� ie �� �e ���  c   ��   f �؅   f �΅  5f    ��a+E ��a�&  ��aT  �b��  �*br�    �u  ]u  l�  �/K  `d;   �o Zo �h  ]�  ��__s �6G  ��$  �Zo ���O  �)G  ��__v �st  ���d�j  �u  ���  %�  �dc   �{o p ���  � ��V  ���  ���  Jf �F�  �d W  ��T�  �f ��d   �o �_�  �f ��  �d   V��  �f   ��d	   �T�  �f ��d	   �_�  	g      ���  ��  e�   �3p �q ��  � ��  ��A�  e8W  �q �O�  g �8W  �Z�  ���  e8W  Ɲ��  g �8W  ���  ���  tg �F�  Se`W  ��T�  �g �Se   �p �_�  �g ��  Xe   V��  h   ��e	   �T�  h ��e	   �_�  (h        �A�  /exW  ��O�  ;h �xW  �Z�  �h ���  /exW  Ɲ��  ;h �xW  ���  �h ���  �h �F�  se�W  ��T�  !i �se   �q �_�  ?i ��  xe   V��  xi   ��e	   �T�  �i ��e	   �_�  �i         ��W   f  �r �w �h  Ӕ  ���|  u�T  ���h  u�T  �� �  u�w ��$r  v�x  ��+�  v�  � �$  w�w �$��*  w�w �(��W  �ȱ  z�w ��w  {�w �i ��  }�w  �i ���  �  j �%  ��  �j �a�  ��t  �j �F�  ��w k �}�  	f   z)s ���  �$ ���  )f�W  �]s �ˆ  hk ���  �k �@f��   �pfq   t �__c �uX  ul �l�  pf   ��s �z�  �l ��  |f   ��s ��   �|f��   �~fc   ���  ��  �l ��  �f   ��.�  m �$�  /m    ��  Pf   �St ��  Bm ���  Vm ���  Pf   ���  Bm ���  jm   ��W  �v ���  ��  m ��  gX  ��t ���  �m �g[e  �0X  �t ��  ��  �m ��  #g   ����  n �1g[e   ���  GgPX  �ru ���  #n ��  QghX  ��,�  ]n �Qg   Ju �7�  �{  Zg   B�+{  �5{  {n   ��h   �,�  �n ��h   �7�      ���  vg   ��u �ˆ  �n ���  �n ��g��   ��X  ��  ��  .o �l�  �g�X  ��z�  no ���  �g�X  ����  no ��X  ���  �o ���  �o �F�  �g�X  ��T�  p ��g   [v �_�  /p ��  �g   V��  Mp   ��h   �T�  `p ��h   �_�  sp         ��X  {w �R'  ��c  ���  h   ��v ���  �p �h�   ��  ,h�X  ��v ���  �p �Ah[e  ���  Ph   �*w �ˆ  �p ���  Hq �`h��   �l�  �hY  �Tw �z�  �q ��h��   ���  �h   ����  ����h�    �fr�    �x  �u  �w  ]u  l�  uX  ��W  i�  ��w ^~ �h  Ӕ  ���|  ��T  ���h  ��T  �� �  �^~ ��$r  ��x  ��+�  ��  � �$  �c~ �$��*  �h~ �(�(Y  �ȱ  �m~ ��w  �r~ �q ��  ��w  
r ���  ��  Vr �V�  �w~ �r �%  ��   s ���  iPY  ��x �ˆ  |s ���  �s �Si��   ��kq   zy �__c �uX  �s �l�  �kpY  �;y �z�   t ��  �k   �0y ��   ��k��   ��Y  �__i ��  9t ��  l   ��.�  dt �$�  wt    �}�  i   ��y ���  �t  ���  �i�Y  ��{ �ˆ  �t ���  �t ���  �i�Y  ԝ�  �t ��  �t �A�  �i�Y  ��z �O�  �t ��Y  �Z�  �t ���  �iZ  ��z ���  �t �Z  ���  �t ���  u �F�  �j8Z  ��T�  zu ��j   �z �_�  �u ��  �j   V��  �u   �k	   �T�  �u �k	   �_�  �u      ���  �iPZ  Ɲ��  �u ���  �v    �A�  �ihZ  ��O�  jw �hZ  �Z�  �w ���  �ihZ  Ɲ��  jw �hZ  ���  �w ���  �w �F�  �j�Z  ��T�  4x ��j   �{ �_�  Rx ��  �j   V��  |x   ��k	   �T�  �x ��k	   �_�  �x          ��Z  �| ���  ��  �x �__c �uX  y �l�  �i�Z  ��| �z�  =y ���  �i�Z  ����  =y ��Z  ���  yy ���  �y �F�  k[  ��T�  z �k   �| �_�  %z ��  k   V��  Cz   ��k	   �T�  Vz ��k	   �_�  iz       �([  �__i ��  |z �@[  �F�  ��w �z    ���  Ojh[  ��} ���  �z ��  Yj�[  ��,�  { �Yj   k} �7�  �{  bj   B�+{  �5{  .{   �Dk   �,�  B{ �Dk   �7�      ��  �j   ��} ��  U{ ���  i{ ���  �j   ���  U{ ���  }{   ���  Cl�[  �~ ���  �{ �Yl�   ��l$   R~ �__i ��  �{ ��  �l�[  ����  �{ ��l[e   �(ir�    �x  �u  �w  ]u  l�  �  ��V  m  ��~ �� �h  Ӕ  ���|  (�T  ���h  (�T  �{ �$  (�� ���*  )�� ��y  )�v  � ��[  �ȱ  ,�� �'y  -�� �{ ��w  .�� �b�  /�� �����  2�j  ����i  3�#  ���}�  m�[  ,w ���  |  �x�  <m@   0� ���  7| ���  |  ���  |m \  1� ���  �D����  �|  �3�  On\  <߁ �[�  �| �O�  �| ���  On\  Ν�  �| ��  �| �A�  On0\  �� �O�  �| �0\  �Z�  �| ���  OnX\  ��� ���  �| �X\  ���  �| ���  } �F�  �nx\  ��T�  g} ��n   ̀ �_�  �} ��  �n   V��  �}   �o	   �T�  S�o	   �_�  P     ���  `n�\  Ɲ��  �} ���  ~    �A�  \n�\  ��O�  f~ ��\  �Z�  �~ ���  \n�\  Ɲ��  f~ ��\  ���  �~ ���  �~ �F�  �n�\  ��T�  �~ ��n   �� �_�    ��n	   �T�   ��n	   �_�            ��  rn
   =.� ��  2 ���  F ���  rn
   ���  2 ���  Z   ��  �n   :}� ��  o ���  � ���  �n   ���  o ���  �   �2m9 �<mr�  �n�w   �u  �w  ]u  3 l�  w�w Ƃ z)l   ��V  0o�  �ނ � �h  Ӕ  ���|  D�T  ���h  D�T  � �$  E� ���*  E� ��y  E�v  � ��\  �ȱ  H� �'y  I�� � ��w  J�� ��  K � ���޲  N�j  ��~��i  O�#  ��~�}�  :o ]  H�� ���  �  � �  bo�   L� ��  	� ��  Q�  ���  �o]  M� ���  ������  d�  �3�  q0]  X)� �[�  w� �O�  �� ���  q0]  Ν�  w� ��  �� �A�  qH]  �g� �O�  �� �H]  �Z�  ǀ ���  qp]  �@� ���  �� �p]  ���  ǀ ���  � �F�  sq�]  ��T�  9� �sq   � �_�  W� ��  xq   V��  u�   ��q	   �T�  S��q	   �_�  P     ���  )q�]  Ɲ��  �� ���  ��    �A�  %q�]  ��O�  8� ��]  �Z�  `� ���  %q�]  Ɲ��  8� ��]  ���  `� ���  �� �F�  �q�]  ��T�  ɂ ��q   �� �_�  ݂  ��q	   �T�  �� ��q	   �_�  ݂          ��  ;q
   Yx� ��  � ���  � ���  ;q
   ���  � ���  ,�   ��  `q   Vǆ ��  A� ���  U� ���  `q   ���  A� ���  i�   �Xo9 �bor�  ��p�w   �u  �w  ]u  3 l�  w�w � z)l   �8X   r=  �(� )� �h  Ӕ  ���|  t�T  ���h  t�T  ��$  t)� ���*  u.� ��y  u�v  � ��l  v�j  �$��]  �ȱ  x3� �'y  y8� ��w  z=� �R'  {�c  ��i  }�#  ���__i ~�  �}�  r
   x	� ���   ��  #r^  {%� ���   ���  Pr0^  � �ˆ  ���  ���  Pr0^  ԰�  ��  �A�  PrX^  �;� �O�  �X^  �Z�  ���  Pr�^  �� ���  ��^  ���  ���  �F�   s�^  ��T�  � s	   �� �T�  � s	   �_�    �t   �_�  ��  t   V��       ���  nr�^  ư��  ���     �A�  cr�^  ��O�  ��^  �Z�  ���  cr�^  ư��  ��^  ���  ���  �F�  `s_  ��T�  �`s   ȉ �_�  ��  is   V��    ��}	   �T�  ��}	   �_�           ���  �r _  �&� ���  ���  ���  � _  �    �@_  y� �__c �q  �XF  ��j  �����  �r�_  ��� ���  ���  ���  ��_  �    ��_  G� ���  ��j  ��  �B� ���Q�  �R� ���Y�  �R� ���ʥ  �b� ���i�  �b� ���|�  �r� ��h  r� ���  	r� ��  �t	   4U� ��  ���  ���  �t	   ���  ���    ��  �u   w� ��  ���   �l�   v   ��� �z�   ���  v�_  �ȋ ���  ���  ���  ��_  �    ��  +v   0� ��  ���  ���  +v   ���  ���    �l�  py   #� �z�   ��_  ٌ �Y�  �j  �����  �y   %`� �ˆ  ���   �l�  3z   &|� �z�   ��  Gz`  &�� ���  ��   �l�  ^z   '�� �z�   ��  rz(`  '���  ��    �l�  @v   ��� �z�   ���  Pv@`  �*� ���  ���  ���  �@`  �    ���  kv5   �F� ���   �l�  0w   �b� �z�   ���  dw   �~� ���   �Ǉ   x   ��� �߇  �Շ   � �  x�   � ��  ��   ���  �x``  �� ���  ���   �x�   y<   �� ���  ���   ���  <yx`  �(� ���  ���   ��  @{   
�'�  ��    ���  ^t�`  ����  ���  ���  ��`  �     �l�  �s�`  :%� �z�  ���  �s�`  ����  ��`  ���  ���  �F�  �t�`  ��T�  ��t   �� �_�  ��  �t   V��    �u	   �T�  �u	   �_�        ��  �s   =d� ��  ���  ���  �s   ���  ���    ���  �t�`  ;� ���  ��  �ta  ��,�  ��t   ȏ �7�  �{  �t   B�+{  �5{    ��~   �,�  ��~   �7�      ��  �s
   B��  ���  ���  �s
   ���  ���      �u  �w  ]u  3 l�  wq  R� z)l  	 w�w b� z)l   w�w r� z)l   w�w �� z)l   �-V  @  ���  � �h  Ӕ  ���|  �T  ~� ��h  �T  Ã �$   � ���*  � ��y  �v  � �0a  �ȱ  	
� �'y  
� � ���  r� �� �}�  W   	N� ���  H�  ��  `   {� �'�  ��  ��  �  �3�  �Ha  �� �[�  �  �O�  �u  ���  �Ha  ΍�  �  ��  �u  �A�  �ha  �ْ �O�  �u  �ha  �Z�  ���  ��a  Ʋ� ���  �u  ��a  ���  ���  g� �F�  ��a  ��T�  �� ��   �� �_�  Մ ��  �   V��  �   �C�	   �T�  V�C�	   �_�  P     ���  ��a  Ɲ��  � ���  ^�    �A�  ��a  ��O�  �� ��a  �Z�  ޅ ���  ��a  Ɲ��  �� ��a  ���  ޅ ���   � �F�  �b  ��T�  G� ��   j� �_�  [�  ��	   �T�  n� ��	   �_�  [�          ��  �   � ��  �� ���  �� ���  �   ���  �� ���  ��   �`9 ���   �u  �w  ]u  3 �mV  `�  �,� �� �h  Ӕ  ���|  �T  �� ��h  �T  � �$  �� ���*  �� ��y  �v  � �(b  �ȱ  �� �'y  �� $� ��h  r� 7� �}�  w�   �� ���  ��  ��  ��   � ��  �}  ���  $�  �3�  ��@b   -� �[�  �  �O�  �  ���  ��@b  ΍�  �  ��  �  �A�  ��`b  �k� �O�  �  �`b  �Z�  ���  ���b  �D� ���  �  ��b  ���  ���  �� �F�  ��b  ��T�  �� ��   � �_�  � ��  �   V��  4�   �c�	   �T�  V�c�	   �_�  P     ���  ʀ�b  Ɲ��  G� ���  ��    �A�  ƀ�b  ��O�  �� ��b  �Z�  � ���  ƀ�b  Ɲ��  �� ��b  ���  � ���  A� �F�  �c  ��T�  �� ��   �� �_�  ��  �'�	   �T�  �� �'�	   �_�  ��          ��  ـ   !|� ��  É ���  ׉ ���  ـ   ���  É ���  �   ���9 ����   �u  �w  ]u  3 A  �� � �h  %~  �__p 	K4  �__c 	Kq  }�%  	N�    ��5  ���  �
� *� Y�  �t  �h  n�  ���|  �O4  ���h  �O4  ��$  �*� ���*  �/� ��#�  �4� � � c  � �e  ��  �k  ��'  ��  ��1  ~ȱ  �9� ��w  �>�  � �ϴ  ��`  �R��k  �ǘ Q� ͘ �� �ԥ  �C� �� ���  ��t  � �x  �l� 8� ��  �u  �� �)�  ��!  �T���  ��j  Ӌ �__n ��j  �� �a�  ��t  8� ��e  ��t  � �/t  ��!  �X�S�  �C� ,� �__p ��'  �\�}�  ��   ��� ���  {�  ���  ǁ   ��� ���  �� �X�  ǁ   	��}�  �p�  �� �f�  (�   ���  �   �D� ���  Ȏ �X�  �   	��}�  �p�  6� �f�  Ȏ   �@c  �� �__i ��j  J� �pc  ���  �t� �� w� ��  ^��c  ;� �3�  �� �'�  � ��  +� ��c  ��  �3�  �'�  ��c  �@�  n� �K�  �V�  �� ��c  �b�  &� �d  �n�  �� �k��e ���f �܈af ��Lf �,�7f      ���  f�(d  g� �ˆ   ���  � ���  f�(d  ԝ�   ��  � �A�  f�Pd  ��� �O�  � �Pd  �Z�  n� ���  f��d  �f� ���  � ��d  ���  n� ���  Ē �F�  ���d  ��T�  !� ���   =� �_�  ?� ��  ��   V��  ]�   �p�   �T�  p� �p�   �_�       ���  ���d  Ɲ��  �� ���  �    �A�  z��d  ��O�  Ԕ ��d  �Z�  � ���  z��d  Ɲ��  Ԕ ��d  ���  � ���  Y� �F�  $� e  ��T�  �� �$�   :� �_�  Օ ��  -�   V��  ��   �@�   �T�  � �@�   �_�           ���  Ђ8e  Ր� ���  %� ����   ���  �Xe  黟 �ˆ  :� ���  \� ���  �Xe  ԝ�  :� ��  \� �A�  ��e  �� �O�  \� ��e  �Z�  ~� ���  ��e  ƺ� ���  \� ��e  ���  ~� ���  ǖ �F�  C�f  ��T�  $� �C�   �� �_�  B� ��  L�   V��  `�   � �   �T�  s� � �   �_�       ���  �(f  Ɲ��  �� ���  ,�    �A�  ��@f  ��O�  �� �@f  �Z�  #� ���  ��@f  Ɲ��  �� �@f  ���  #� ���  l� �F�  ��f  ��T�  �� ��   �� �_�  ܙ ��  ��   V��  �   �0�   �T�  � �0�   �_�           ��f  Ǣ �__c ��5  ,� �__q �C� �l�  ��f  묠 �z�  `� ���  ��f  ����  `� ��f  ���  �� ���  ؚ �F�  ���f  ��T�  � ���   �� �_�  ;� ��  ��   V��  Y�   �`�   �T�  l� �`�   �_�        �I  5�   �� �m  � �`  Ǜ �S  �� �C�Bg  ���  [�g  � �Ȍ  7� ���  `� ���  [�g  	���  7� ��  `� �g  ��  �� �Mz  [�   	/�� �[z  `� �4z  [�   	��Bz  `� �z  [�   	-�$z  `�    ��~  ��   	2ȡ ��~  �� ��~  Ȝ  �4z  ��   	3� �Bz  �� �z  ��   	-�$z  ��   �  �� g  	3�� �#  � �   � ���    �#  B� �  U� ��{  ��   	�f� ��{   ��~  ��   	װ�~  ��~  j�    �}�3     ���  ��   �Ȍ  �� ���  �� �
���    ���  ��8g  �^� ���  Ý ��  ��Xg  ��,�  � ���   6� �7�  �{  ��   B�+{  �5{  �   ���#   �,�  � ���#   �7�      �֌  �   �� ��  *� �Mz  �   	6�[z  *�   �pg  �� �R'  Ŵ� ?� l� �__j �l� ^� ���  ���g  ��� �ˆ  }� ���  �� ���  ���g  ԝ�  }� ��  �� �A�  ���g  �� �O�  �� ��g  �Z�  �� ���  ���g  �� ���  �� ��g  ���  �� ���  �� �F�  0� h  ��T�  � �0�   �� �T�  ,� �0�   �_�    ���   �_�  ?� ��  ��   V��  ]�      ���  Ɋh  Ɲ��  p� ���  ��    �A�  0h  ��O�  :� �0h  �Z�  \� ���  0h  Ɲ��  :� �0h  ���  \� ���  �� �F�  c�`h  ��T�  Р �c�   ǥ �_�  � ��  l�   V��  �   � �   �T�  +� � �   �_�           �l�  �xh  �� �z�  >� �����   ���  ���h  ǝ��  x� ��  ���h  ��,�  �� ���   �� �7�  �{  ��   B�+{  �5{  ��   ���    �,�  �� ���    �7�       ���   �   � �ˆ  ҡ ���  $� �0���   �l�  ���h  �� �z�  ^� ���  ���h  ����  ^� ��h  ���  �� ���  �� �F�  Ɔ�h  ��T�  � �Ɔ   �� �_�  5� ��  φ   V��  S�   �0�   �T�  f� �0�   �_�        ���  ���h  I� ���  y� ��  �i  ��,�  �� ��   !� �7�  �{  �   B�+{  �5{  ƣ   ��   �,�  ڣ ��   �7�      �l�  V�   s� �z�  � �b���   ���  ~�'   �� ���  � ����   ���  ��   �Ш �ˆ  /� ���  �� �����   ���  ،0i  ��� ���  �� ����   ���  �   �,� �ˆ  Ф ���  "� �����   �l�  F�Hi  �U� �z�  \� �R���   �l�  W�`i  �~� �z�  �� �c���   �s��    ��  6�   Q٩ ��  �� ���  ʥ ���  6�   ���  �� ���  ޥ   �3�  <�   V� �[�  � �O�  I� �F���   ��  \�xi  ��� ���  �� �4z  \��i  	#K� �Bz  ��  ��}  e��i  	#��}  � ��}  1� ����  �Ru[   ��  p��i  X�� ���  O� �4z  p�   	#ê �Bz  O�  ��}  v��i  	#��}  �� ��}  ǧ �Ԏ��  �Ru`   ��i  � �gh  %C� � �__i 'l� � ���  ��j  (\� �ˆ  E� ���  Z� ����   �l�  �(j  )�� �z�  o� ����   ���  '�@j  (���  �� ��  1�Xj  ��,�  �� �1�   � �7�  �{  6�   B�+{  �5{  ��   �I�   �,�  ˨ �I�   �7�       �Mz  p�   2;� �[z  ި  �y�7   �� �z  4�� � ��x  5u  +� �Mz  ��   7�� �[z  C�  ����  ����!  ��  ��    ;L� ��  X� ���  x� �~  ��pj  	\/� �~  x� �4z  ��   	<$� �Bz  x� �z  ��   	-�$z  x�   �Ѕ�	   �z  Ѕ   	]�$z  ʩ   ��  ۅ   <�� �#�  � �~  ۅ   	h�~  � ���	    ��� �!   <� �˗ 1� ��� ��� F� ��!   �ٗ s� �fz  ��j  	P�� �tz  ��  ��h    �Mz  �   ?!� �[z  ��  ���  )��j  BU� �Ȍ  Ԫ ���  3� �9���   ��  ��   G�� ��  Q� ���  e� ���  ��   ���  Q� ���  y�   ��  ��   W� ��  �� ���  �� ���  ��   ���  �� ���  ��   ��  �   �j� ���  ˫ �4z  �   	#1� �Bz  ˫  ��}  ��   	#��}  � ��}  � �	���  �Ru[   ��  	�   X� ���  u\��4z  	�   	#�� �Bz  u\� ��}  �   	#��}   � ��}  M� ����  �Ru`   ���r�  ���M! ��3  ���3  �K�j  �}�A   �'�Ge  �u  �w  �x  ]u  l�  �5  ��5  0��  �k� �� Y�  �t   �h  n�  ���|  �O4  ���h  �O4  ��$  ��� ���*  ��� ��#�  ��� � ��j  �� �e  ��  �k  ��'  ��  �B,  ~ȱ  ��� ��w  ��� `� �ϴ  �,a  �R��k  �(� �� .� � �ԥ  �C�  � ���  ��t  l� �x  �Ͱ �� ��  �u  � �)�  ��!  �T���  ��j  3� �__n ��j  _� �a�  ��t  �� ��e  ��t  l� �/t  ��!  �X�S�  �C� �� �__p ��'  �\�}�  9�   �� ���  ۯ  ���  w�   �Z� ���  �� �X�  w�   	��}�  �p�  \� �f�  ��   ���  ��   ��� ���  (� �X�  ��   	��}�  �p�  �� �f�  (�   ��j  �� �__i ��j  �� �k  ���  �ղ � ذ ��  �Hk  �� �3�  � �'�  O� ��  �� �hk  ��  �3�  �'�  �hk  �@�  β �K�  �V�  � ��k  �b�  �� ��k  �n�  � ���e �j�f ���af ���Lf �ܖ7f      ���  ��k  ȵ �ˆ  "� ���  x� ���  ��k  ԝ�  "� ��  x� �A�  ��k  �� �O�  x� ��k  �Z�  δ ���  �(l  �Ǵ ���  x� �(l  ���  δ ���  $� �F�  C�Pl  ��T�  �� �C�   �� �_�  �� ��  L�   V��  ��   � �   �T�  е � �   �_�       ���  5�hl  Ɲ��  � ���  |�    �A�  *��l  ��O�  4� ��l  �Z�  c� ���  *��l  Ɲ��  4� ��l  ���  c� ���  �� �F�  Ԕ�l  ��T�  � �Ԕ   �� �_�  5� ��  ݔ   V��  _�   ��   �T�  r� ��   �_�           ���  ���l  �� ���  �� �0��   ���  ���l  �� �ˆ  �� ���  �� ���  ���l  ԝ�  �� ��  �� �A�  ��0m  �B� �O�  �� �0m  �Z�  ޸ ���  ��xm  �� ���  �� �xm  ���  ޸ ���  '� �F�  ��m  ��T�  �� ��   � �_�  �� ��  ��   V��  ��   ���   �T�  ӹ ���   �_�       ���  ���m  Ɲ��  � ���  ��    �A�  ���m  ��O�  T� ��m  �Z�  �� ���  ���m  Ɲ��  T� ��m  ���  �� ���  ̻ �F�  ��(n  ��T�  � ���   � �_�  <� ��  ��   V��  f�   ���   �T�  y� ���   �_�           �@n  (� �__c ��5  �� �__q �C� �l�  ɐpn  �� �z�  �� ���  ɐpn  ����  �� �pn  ���  	� ���  8� �F�  3��n  ��T�  }� �3�   � �_�  �� ��  <�   V��  ��   ��   �T�  ̽ ��   �_�        �I  �   �J� �m  ߽ �`  '� �S  _� ��Bg  ���  ��n  ��� �Ȍ  �� ���  �� ���  ��n  	���  �� ��  �� ��n  ��  � �Mz  �   	/�� �[z  �� �4z  �   	��Bz  �� �z  �   	-�$z  ��    ��~  6�   	2)� ��~   � ��~  (�  �4z  ;�   	3e� �Bz  @� �z  ;�   	-�$z  @�   �  >��n  	3� �#  b� �  �� �P�    �#  �� �  �� ��{  P�   	�Ǻ ��{   ��~  Z�   	װ�~  ��~  ʿ    �-�3     ���  ��   �Ȍ  � ���  �� �����    ���  L��n  鿻 ���  #� ��  V��n  ��,�  E� �V�   �� �7�  �{  _�   B�+{  �5{  c�   �p�#   �,�  w� �p�#   �7�      �֌  đ   �� ��  �� �Mz  đ   	6�[z  ��   �o  � �R'  �� �� Ͱ �__j �Ͱ �� ���  `�(o  �U� �ˆ  �� ���  �� ���  `�(o  ԝ�  �� ��  �� �A�  `�Po  �{� �O�  �� �Po  �Z�  � ���  `��o  �T� ���  �� ��o  ���  � ���  � �F�  ���o  ��T�  n� ���    � �T�  �� ���   �_�    �C�   �_�  �� ��  H�   V��  ��      ���  y��o  Ɲ��  �� ���  �    �A�  r��o  ��O�  �� ��o  �Z�  �� ���  r��o  Ɲ��  �� ��o  ���  �� ���  �� �F�  � p  ��T�  0� ��   (� �_�  N� ��  �   V��  x�   ���   �T�  �� ���   �_�           �l�  ��p  �~� �z�  �� �����   ���  `�0p  ǝ��  �� ��  j�Hp  ��,�  �� �j�   � �7�  �{  o�   B�+{  �5{  �   ���    �,�  � ���    �7�       ���  В   F� �ˆ  2� ���  �� �����   �l�  `�`p  � �z�  �� ���  `�`p  ����  �� �`p  ���  �� ���  � �F�  v��p  ��T�  w� �v�   � �_�  �� ��  �   V��  ��   ���   �T�  �� ���   �_�        ���  ���p  �� ���  �� ��  ���p  ��,�  � ���   �� �7�  �{  ��   B�+{  �5{  &�   �͚   �,�  :� �͚   �7�      �l�  �   �� �z�  M� ����   ���  .�'   �� ���  z� �B��   ���  U�   �1� �ˆ  �� ���  �� �e���   ���  ���p  �Z� ���  � �A��   ���  ��   ׍� �ˆ  0� ���  �� �����   �l�  ���p  Ҷ� �z�  �� ����   �l�  � q  ��� �z�  �� ����   �#��    ��  �   Q:� ��  � ���  *� ���  �   ���  � ���  >�   �3�  �   Vn� �[�  S� �O�  �� �����   ��  �q  ��� ���  �� �4z  �8q  	#�� �Bz  ��  ��}  �Pq  	#��}  H� ��}  �� �����  �Ru[   ��   �hq  X]� ���  �� �4z   �   	#$� �Bz  ��  ��}  &��q  	#��}  �� ��}  '� �����  �Ru`   ��q  |� �gh  %C� e� �__i 'Ͱ y� ���  ���q  (�� �ˆ  �� ���  �� �����   �l�  ���q  )�� �z�  �� �ɛ��   ���  כ�q  (���  �� ��  ��q  ��,�  �� ��   S� �7�  �{  �   B�+{  �5{  �   ���   �,�  +� ���   �7�       �Mz   �   2�� �[z  >�  �)�7   � �z  4� x� ��x  5u  �� �Mz  E�   7�� �[z  ��  �9��  �]��!  ��  f�    ;�� ��  �� ���  �� �~  f�r  	\�� �~  �� �4z  f�   	<�� �Bz  �� �z  f�   	-�$z  ��   ����	   �z  ��   	]�$z  *�   ��  ��   <�� �#�  d� �~  ��   	h�~  d� ����	    ��� ��!   <b� �˗ �� ��� ��� �� ���!   �ٗ �� �fz  ��(r  	PV� �tz  ��  ���h    �Mz     ?�� �[z  ��  ���  ٓ@r  B�� �Ȍ  4� ���  �� ����   ��  c�   G� ��  �� ���  �� ���  c�   ���  �� ���  ��   ��  C�   WT� ��  �� ���  � ���  C�   ���  �� ���  �   ��  ��   ��� ���  +� �4z  ��   	#�� �Bz  +�  ��}  ��   	#��}  @� ��}  m� �����  �Ru[   ��  ��   XC� ���  u\��4z  ��   	#
� �Bz  u\� ��}  ��   	#��}  �� ��}  �� �Μ��  �Ru`   �E�r�  �T��. ���3  ���3  ���j  �-�A   �לGe  �u  �w  �x  ]u  l�  � 5  ���   ��� F� �h  n�  ���|  mO4  �� ��h  mO4  ����  m�t  ��$  mF� ���*  nK� � �#�  nP� �$�`r  ;� ��^  p�!  �X���  ��   p�� ���  � �X�  ��   	��}�  �p�  \� �f�  �   ��  D��r  t�� ���  �� ��}  D��r  	#a� ��}  �� ��}  �� ���   ��}  � ��}  "� �q}  ���r  	�U� ��}  5� �{}  J� ��y  ���r  
V��y  5� ��y  J� ��r  �	z  _�    ����    �4z  L�   	#�Bz  �� �z  L�   	-�$z  ��    ��  ��   t� ���  u`��4z  ��   	#�� �Bz  u`� ��}  ��   	#��}  r� ��}  �� �Ý��  �Rud   ��� �,�T  �A�5j  ���I�  �̝Ge  �u  �w  x  �e5  Н�  �m� � �h  n�  ���|  zO4  �� ��h  zO4  ����  z�t  ��$  z� ���*  {
� � �{�  {� �$��r  �� T�e  }�  �ȱ  � ��w  �� �� ��^  ��!  �\�R'  �0� � �� �}�  ٝ s  U� ���  <�  ���  �   ��� ���  \� �X�  �   	��}�  �p�  �� �f�  \�   �Mz  )�s  ��� �[z  �� �4z  )�   	��Bz  �� �z  )�   	-�$z  ��    ��  <�0s  ��� ���  �� �4z  <�   	#8� �Bz  ��  ��}  B�Xs  	#��}  -� ��}  \� ��0   ��}  z� ��}  �� �q}  �xs  	��� ��}  �� �{}  �� ��y  �xs  
V��y  �� ��y  �� �xs  �	z  ��    �.��     �.�  ���s  �� �F�  � �<�  "� ����   ��  ���s  ��� ��  6� ���  �~  ���s  	\�~  �4z  ���s  	<�� �Bz  �z  ���s  	-�$z    ����	    �T�  Ğ   ��� �b�  V� �z  Ğ   	&�$z  V�   ���  ʞ�s  �c� �Ʊ  x� ���  �� ���  3� ���  �� �!�  �   �X� �S�  �� �F�  �� �9�  �� �/�  �� ��#e  �	��c   ��  X�   ��� ���  ud��4z  X�   	#�� �Bz  ud� ��}  ^�   	#��}  �� ��}   � �m���  �Ruc   ��r�  ��� ���I�  �v�Ge  �u  �w  	x  ]u  l�  �8B  ���
  �6� Y� �h  ��  ���|  �D6  ���h  �D6  ��$  �Y� ���*  �^� ����  �c� � ��s  N� ��  ��=  �ϴ  �ia  �Z~ȱ  �h� ��k  ��� 3� �� �� �ԥ  ��j  g� �__c �y?  �� � �  ��t  � ���  ��t  �� ���  ��j  �� ��  ˧t  �� �L}  ̧t  f� �p�  ��!  �\�S�  �m� v� �}�  ��   ��� ���  ��  �3�  �� t  ��� �[�  
� �O�  �� �����   �8t  �� �r  �u  �� �l�   �Xt  ��� �z�  � ����   ���  �pt  �/� �Ȍ  n� ���  �� �1���   ���  1�   �X� ���  �� �D��   ���  N�   ��� �ˆ  �� ���  �� �^���   �l�  i�   ��z�  4� �u���    ���  ���t  ��� �ˆ  a� ���  �� ���  ���t  ԝ�  a� ��  �� �A�  ���t  ��� �O�  �� ��t  �Z�  �� ���  ���t  Ɲ��  �� ��t  ���  �� ���  � �F�  ��u  ��T�  U� ���   �� �_�  s� ��  ��   V��  ��   ���   �T�  �� ���   �_�  ��        �A�  �� u  ��O�  �� � u  �Z�  �� ���  ��Xu  Ʒ� ���  �� �Xu  ���  �� ���  �� �F�  ���u  ��T�  =� ��u  �� �_�  [� ��  ��   V��  y�   �`�	   �T�  �� �`�	   �_�  ��      ���  ���u  Ɲ��  �� ���  �      ���  ҟ�u  �+� ���  �� �X�  ҟ�u  	��}�  �p�  �� �f�  ��   ��u  r� ~9�  ��t  �:�   �   ֒� �m�  �� �`�  "� �[�  f� �Q�  �� � �   �{�  ��   ���  �   ��� �Ȍ  J� ���  ]� ����   ���  ��v  ��� �Ȍ  }� ���  �� ����   ���  �(v  �� ���  �� ��  �Hv  ��,�  /� �hv  c� �7�  �{  %��v  B�+{  �5{  M�   �0�   �,�  a� �0�   �7�      ���  5��v  �� �ˆ  t� ���  �� ���  5��v  ԝ�  t� ��  �� �A�  5��v  ��� �O�  �� ��v  �Z�  �� ���  5� w  Ƶ� ���  �� � w  ���  �� ���  � �F�  5�(w  ��T�  S� �5�   �� �_�  q� ��  >�   V��  ��   ���   �T�  �� ���   �_�       ���  K�@w  Ɲ��  �� ���  �    �A�  A�Xw  ��O�  �� �Xw  �Z�  �� ���  A�Xw  Ɲ��  �� �Xw  ���  �� ���  �� �F�  ��w  ��T�  H� ��   �� �_�  f� ��  �   V��  ��   ��   �T�  �� ��   �_�           ��w  D� �r  �u  �� �l�  a��w  �� �z�  � ��  s�   �	� ��   �m���   ���  ���w  �Ȍ  T� ���  g� �����    ���  @�   �w� �Ȍ  �� ���  �� �M���   ���  "� x  �
� ���  �� ��  0�(x  ��,�  �� �Hx  �� �7�  �{  9�`x  B�+{  �5{  ��   �`�   �,�  � �`�   �7�      ���  I�xx  �1� �ˆ  #� ���  E� ���  I�xx  ԝ�  #� ��  E� �A�  I��x  �W� �O�  E� ��x  �Z�  g� ���  I��x  �0� ���  E� ��x  ���  g� ���  �� �F�  I��x  ��T�  �� �y  � �_�  �� ��  R�   V��  "�   ���   �T�  5� ���   �_�       ���  c� y  Ɲ��  H� ���  ��    �A�  U�8y  ��O�  � �8y  �Z�  4� ���  U�8y  Ɲ��  � �8y  ���  4� ���  c� �F�  ϡpy  ��T�  �� �ϡ   � �_�  �� ��  ء   V��  ��   ���   �T�  � ���   �_�           �l�  �   ��z�  � ��  ��   �f� ��   �����    ��y  �� �__q .m� �I  2�   /�� �m  C� �`  �� �S  �� �C�Bg  ���  Q��y  2�� �Ȍ  � ���  � �c���   ���  ��   </� �Ȍ  ?� ���  S� �
���   ���  ��y  =c� �Ȍ  �� ���  �� ����   ���  ��y  A�� ���  �� ��  '�z  ��,�  �� �'�   �� �7�  �{  0�   B�+{  �5{  �   �Щ    �,�  0� �Щ    �7�      ���  =�   A/� �ˆ  C� ���  �� �M���   � z  �r  Du  � �l�  X�@z  C�� �z�  *� ��  j�   ��� ��   �d���   ���  ��Xz  I�Ȍ  q� ���  �� �����     �Mz  ��   $�� �[z  ��  ���  ��   %� �Ȍ  �� ���  �� �����   ���  ��   &E� �Ȍ  � ���  '� �����   ���  �pz  y� �Ȍ  G� ���  ~� ����   ��  +�    �� ��  �� �Mz  +��z  	.�� �[z  ��  �?��	   ���  o��z  WW� ���  �� ��  }��z  ��,�  �� ��z  /� �7�  �{  �� {  B�+{  �5{  �   �Х   �,�  � �Х   �7�      ���  ��{  W� �ˆ  2� ���  T� ���  ��{  ԝ�  2� ��  T� �A�  ��@{  ��� �O�  T� �@{  �Z�  v� ���  ��p{  �~� ���  T� �p{  ���  v� ���  �� �F�  ���{  ��T�  �� ��{  U� �_�  � ��  ��   V��  1�   � �   �T�  D� � �   �_�       ���  ���{  Ɲ��  W� ���  ��    �A�  ���{  ��O�  � ��{  �Z�  3� ���  ���{  Ɲ��  � ��{  ���  3� ���  b� �F�  N�|  ��T�  �� �N�   R� �_�  �� ��  W�   V��  ��   �`�   �T�  � �`�   �_�           �l�  £   X�� �z�  !� ��  Σ   ��� ��   �Σ��   �Mz  y�(|  _� �[z  N� �4z  y�H|  	��Bz  N� �z  y�h|  	-�$z  N�    ��  ���|  k�� ���  �� �4z  ��   	#[� �Bz  ��  ��}  ���|  	#��}  �� ��}  � ����  �Ruc   ���  f��|  �'� ���  C� ��  x��|  ��,�  e� �}  �� �7�  �{  ��0}  B�+{  �5{  ��   �0�   �,�  �� �0�   �7�      ���  ��#   c[� �Ȍ  �� ���  �� �����   �l�  ̨   � �z�  �� �ب��   ���  �H}  ��� �Ȍ  � ���  +� �����   ��  W�   k/� ���  ud��4z  W�   	#�� �Bz  ud� ��}  ]�   	#��}  K� ��}  x� �l���  �Ruc   ���+E ���j  ��3   �u�Ge  �u  �w  �x  ]u  bE  �/D  ��k  ��� e� �h  ��  ���|  ��?  �� ��h  ��?  �� �$  �e� ���*  �j� ��__v �o� � �`}  Z� ���  ��!  �X���  ��
   �P� ���  �� �X�  ��
   	��}�  �p�  � �f�  ��   �3�  ��}  �`� �[�  1� �O�  I� ���  ��}  Ν�  1� ��  I� �A�  ��}  ��� �O�  I� ��}  �Z�  a� ���  ��}  �{� ���  I� ��}  ���  a� ���  v� �F�  C��}  ��T�  �� �C�   R� �_�  �� ��  H�   V��  �   �`�   �T�  /� �`�   �_�       ���   �~  Ɲ��  N� ���  ��    �A�  �� ~  ��O�  � � ~  �Z�  F� ���  �� ~  Ɲ��  � � ~  ���  F� ���  u� �F�  P�P~  ��T�  �� �P�   3� �_�  ��  ���   �T�  �� ���   �_�           ��  �   ��� ��  � ���  � ���  �   ���  � ���  +�   ��  !�h~  ��� ���  @� �4z  !��~  	#
� �Bz  @� �z  !�   	-�$z  @�   ��}  *��~  	#��}  o� ��}  �� ���    ��}  �� ��}  �� �q}  ���~  	��� ��}  �� �{}  �� ��y  ���~  
V��y  �� ��y  �� ��~  �	z  �    ����     ��  ͫ   �1� ���  u`��4z  ͫ   	#�� �Bz  u`� ��}  ӫ   	#��}  .� ��}  [� ����  �Rud   ���3  ���� �ӪT  ��Yj   ��Ge  �u  �w  �x  �oD  �k  ��� f� �h  ��  ���|  ��?  n� ��h  ��?  �� �$  �f� ���*  �k� ��__v �p� � ��~  [� ���  ��!  �X���  ��
   �Q� ���  �� �X�  ��
   	��}�  �p�   � �f�  ��   �3�  X��~  �a� �[�  � �O�  ,� ���  X��~  Ν�  � ��  ,� �A�  X�  ��� �O�  ,� �  �Z�  D� ���  X�@  �|� ���  ,� �@  ���  D� ���  Y� �F�  ��`  ��T�  �� ���   S� �_�  �� ��  ��   V��  ��   �Ь   �T�  � �Ь   �_�       ���  p�x  Ɲ��  1� ���  ��    �A�  l��  ��O�  �� ��  �Z�  )� ���  l��  Ɲ��  �� ��  ���  )� ���  X� �F�  ���  ��T�  �� ���   4� �_�  ��  � �   �T�  �� � �   �_�           ��  ��   ��� ��  �� ���  �� ���  ��   ���  �� ���  �   ��  ���  ��� ���  #� �4z  ���  	#� �Bz  #� �z  ��   	-�$z  #�   ��}  ���  	#��}  R� ��}  �� � �    ��}  �� ��}  �� �q}   �(�  	��� ��}  �� �{}  �� ��y   �(�  
V��y  �� ��y  �� �(�  �	z  ��    ���     ��  =�   �2� ���  u`��4z  =�   	#�� �Bz  u`� ��}  C�   	#��}    ��}  >  �R���  �Rud   ��3  �/�� �C�T  �X�}j   �[�Ge  �u  �w  �x  ��D  `�k  ��� g� �h  ��  ���|  ��?  Q  ��h  ��?  �  �$  �g� ���*  �l� ��__v �q� � �@�  \� ���  ��!  �X���  l�
   �R� ���  �  �X�  l�
   	��}�  �p�  �  �f�  �    �3�  ȭ`�  �b� �[�  �  �O�   ���  ȭ`�  Ν�  �  ��   �A�  ȭ��  ��� �O�   ���  �Z�  ' ���  ȭ��  �}� ���   ���  ���  ' ���  < �F�  #�Ѐ  ��T�  � �#�   T� �_�  � ��  (�   V��  �   �@�   �T�  � �@�   �_�       ���  ��  Ɲ��   ���  l    �A�  ܭ �  ��O�  � � �  �Z�   ���  ܭ �  Ɲ��  � � �  ���   ���  ; �F�  0�0�  ��T�  � �0�   5� �_�  �  ���   �T�  � ���   �_�           ��  �   ��� ��  � ���  � ���  �   ���  � ���  �   ��  �H�  ��� ���   �4z  �h�  	#� �Bz   �z  �   	-�$z     ��}  
���  	#��}  5 ��}  d �p�    ��}  � ��}  � �q}  p���  	��� ��}  � �{}  � ��y  p���  
V��y  � ��y  � ���  �	z  �    ����     ��  ��   �3� ���  u`��4z  ��   	#�� �Bz  u`� ��}  ��   	#��}  � ��}  ! �®��  �Rud   �~�3  ���� ���T  �ȭ5j   �ˮGe  �u  �w  x  �gE  Ю�  ��� 0 ]T  %   �h  ��  ���|  rD6  ���h  rD6  ��$  r0 ���*  s5 ��__v s: � ���  % Tߠ  w�l  T��  x�=  �ϴ  yia  �Z�ȱ  z? ��k  {D� 4 J� 
� �ԥ  |�j  � �__c }y?  = ��m  ��$  �'�  �u   ���  ��j  � � �  ��t  � ���  ��t  � �Qr  ��t  $	 ���  ��j  �	 �R'  ��c  �
 �p�  ��!  �\���  ��t   ���  ��t  i ��  �8� � �� �ڪ  �8� D ��T  ��� � �9�  ��j  3 �S�  �m� i �}�  ܮ   z�� ���  8  �(�  �Ё  ��� �>�  J�2�  z  �3�  ��  ��� �[�  � �O�  e �$���   �l�  2� �  �A� �z�  � ��  D�   �6� ��   �>���   ���  o�   �k� ���  ? ���   ���  ��   ��� �ˆ  a ���  � �����   ���  ̯   ��� ���  � �X�  ̯   	��}�  �p�  - �f�  �   �:�  ��  �~� �m�  M �`�  m �[�  � �Q�  � ��&   A� �{�  �  �8�  �Q�  M �[�  m �`�  � �m�  �8�  �{�  �    ���  J�X�  �� ���  � ��  ]���  ��,�    ���  �� �7�  �{  f���  B�+{  �5{     ���   �,�  2 ���   �7�      ���  v�Ђ  �:� �ˆ  E ���  g ���  v�Ђ  ԝ�  E ��  g �A�  v���  �`� �O�  g ���  �Z�  � ���  v�(�  �9� ���  g �(�  ���  � ���  � �F�  v�H�  ��T�  � �`�  � �_�   ��  �   V��  D   ���   �T�  W ���   �_�       ���  ��x�  Ɲ��  j ���  �    �A�  ����  ��O�  � ���  �Z�  � ���  ����  Ɲ��  � ���  ���  � ���  � �F�  ,�ȃ  ��T�  1 �,�   � �_�  O ��  5�   V��  y   � �   �T�  � � �   �_�           �l�   �   � �z�  � ��  /�   �t� ��   �,���   ���  �� �__q 
m� �I  P�   �m  � �`  � �S   �`�Bg   ���  ;�   �� �Ȍ  6 ���  m �K���   ���  ����  �� ���  � ��  �� �  ��,�  � �@�  q� �7�  �{  ��X�  B�+{  �5{  �   �`�   �,�  � �`�   �7�      ���  ��p�  �� �ˆ   ���  # ���  ��p�  ԝ�   ��  # �A�  ����  ��� �O�  # ���  �Z�  E ���  ��Ȅ  ��� ���  # �Ȅ  ���  E ���  g �F�  ���  ��T�  � � �  �� �_�  � ��  ��   V��      ���   �T�   ���   �_�       ���  γ�  Ɲ��  & ���  x    �A�  ��0�  ��O�  � �0�  �Z�   ���  ��0�  Ɲ��  � �0�  ���   ���  N �F�  �h�  ��T�  � ��   �� �_�  � ��  �   V��  �   �P�   �T�  � �P�   �_�           �l�  E���  ��� �z�   ���  E���  ����   ���  ���  / ���  Q �F�  _���  ��T�  � �_�   c� �_�  � ��  h�   V��  �   ��   �T�  � ��   �_�        �Mz  ��   %�� �[z  � �4z  ��   	��Bz  � �z  ��   	-�$z  �    ��  ߰   E4  ��  A ���  U ���  ߰   ���  A ���  i   ��  ���  F�  ���  ~ �4z  �   	#s  �Bz  ~  ��}  �؅  	#��}  � ��}  � �#���  �Ruc   ���  ���  (�  �Ȍ   ���  ( �!���   �Mz  Q�   28 �[z  � �4z  Q�   	��Bz  � �z  Q�   	-�$z  �    �l�  ��   �} �z�  � ��  ��   �r ��   �����   ���  *��  � ���  � ��  4�(�  ��,�   �4�   � �7�  �{  =�   B�+{  �5{      ��+   �,�  4 ��+   �7�      ���  J�   �I �ˆ  G ���  v �W���   �l�  ��@�  �� �z�  � ��  Ӷ   �� ��   �̶��   ��  ��   F ���  ud��4z  ��   	#� �Bz  ud� ��}  ��   	#��}  � ��}  $ �����  �Ruc   ��+E �6�j  ���3   ���Ge  �u  �w  }x  ]u  �B  R � �h  ��  ��|  ��?  ��h  ��?  �$  �� ��*  �� �__v ��  �u  �w  }x  �D q�  ��7   �� 
 �R ��\ ��i ��v ��� ��� � �ηv�  ��?  �|   �" � �h  ��  ��e  ��?  ���h  ��?  ��$  �� ���*  �� ��__v �� � �D ��&   ��� 7 �� K �v _ �i �\ �R ~ � �v�   �u  �w  }x  �oB  `�d  �� �
 �h  ��  ���|  N�?  ���h  N�?  ��$  N�
 ���*  O�
 ��__v O�
 � �X�  � �__l V%   �\�3�  ̸p�  `� �[�  �O�  ����   ��  ��   a� ��  � ���  � ���  ��   ���  � ���  �   ���v�  ���  T��  g�=  �ϴ  hia  �\�ȱ  i�
 ��k  j4 � : � �<�  l�t  q  �+�  m�t  ! �\�  n�t  ~! ��  o�t  �! � �  p�t  " �__n q�  �" �}�  �   i� ���  �"  ���  y
 �__c zbE  # �3�  ]�І  t	 �[�  ## �O�  y# ���  ]�І  Ν�  ## ��  y# �A�  ]� �  �6 �O�  y# � �  �Z�  �# ���  ]�0�  � ���  y# �0�  ���  �# ���  %$ �F�  �P�  ��T�  �$ ��   � �_�  �$ ��  ��   V��  �$   �8�	   �T�  �$ �8�	   �_�  	%      ���  ��h�  Ɲ��  % ���  �%    �A�  t���  ��O�  �& ���  �Z�  ' ���  t���  Ɲ��  �& ���  ���  ' ���  z' �F�  ����  ��T�  �' ���   � �_�  �' ��  ��   V��  !(   �h�	   �T�  4( �h�	   �_�  G(          �l�  ��Ї  z�	 �z�  Z( ���  ��Ї  ����  Z( �Ї  ���  �( ���  ) �F�  ���  ��T�  X) ��   �	 �_�  v) ��  �   V��  �)   ���	   �T�  �) ���	   �_�  �)       ���  ���  ����  �) ��  �(�  ��,�  �) ��   P
 �7�  �{  �   B�+{  �5{  *   ��   �,�  !* ��   �7�       ��  ��   ��
 ��  4* ���  H*  �&�+E   �u  �w  wx  ]u  ��E  м�  ��
 } ]T  �j  �h  ��  ���|  rD6  ���h  rD6  ��$  r} ���*  s� ��__v s� � �@�  r Tߠ  w2s  T��  x�=  �ϴ  yia  �Z�ȱ  z� ��k  {� \* � W �ԥ  |�j  �* �__c }y?  e+ ��m  ��$  �'�  �u  B, ���  ��j  �, � �  ��t  �, ���  ��t  . �Qr  ��t  i. ���  ��j  �. �R'  ��c  �/ �p�  ��!  �\���  ��t  W0 ���  ��t  �0 ��  �� U1 K �ڪ  �� �1 ��T  �K h2 �9�  ��j  �2 �S�  �m� D3 �}�  ܼ   z� ���  4  �(�  �`�  � �>�  J�2�  P4  �3�  �x�  �I �[�  o4 �O�  ;5 �$���   �l�  2���  �� �z�  �5 ��  D�   �� ��   �>���   ���  o�   �� ���  6 ���   ���  ��   �� �ˆ  76 ���  Y6 �����   ���  ̽   �8 ���  �6 �X�  ̽   	��}�  �p�  7 �f�  �6   �:�  ���  �� �m�  #7 �`�  C7 �[�  o7 �Q�  �7 ��&   � �{�  �7  �Ȉ  �Q�  #8 �[�  C8 �`�  k8 �m�  �Ȉ  �{�  �8    ���  B��  �_ ���  �8 ��  U��  ��,�  �8 �0�  7 �7�  �{  ^�H�  B�+{  �5{  �8   �p�   �,�  9 �p�   �7�      ���  n�`�  �� �ˆ  9 ���  =9 ���  n�`�  ԝ�  9 ��  =9 �A�  n���  �� �O�  =9 ���  �Z�  _9 ���  n���  Ɔ ���  =9 ���  ���  _9 ���  �9 �F�  n�؉  ��T�  �9 ���  ] �_�  �9 ��  w�   V��  :   ���   �T�  -: ���   �_�       ���  ���  Ɲ��  @: ���  �:    �A�  z� �  ��O�  d; � �  �Z�  �; ���  z� �  Ɲ��  d; � �  ���  �; ���  �; �F�  �X�  ��T�  < ��   Z �_�  %< ��  �   V��  O<   ���   �T�  b< ���   �_�           �l�   �   � �z�  u< ��  �   �� ��   ����   �p�   �__q 
m� �I  0�   �m  �< �`  �< �S  �< �@�Bg   ���  �   �R �Ȍ  
= ���  A= �+���   ���  x���  � ���  n= ��  ����  ��,�  �= �Њ  � �7�  �{  ���  B�+{  �5{  �=   �@�   �,�  �= �@�   �7�      ���  �� �   �ˆ  �= ���  �= ���  �� �  ԝ�  �= ��  �= �A�  ��(�  �4 �O�  �= �(�  �Z�  > ���  ��X�  � ���  �= �X�  ���  > ���  ;> �F�  ��x�  ��T�  �> ���  � �_�  �> ��  ��   V��  �>   �p�   �T�  �> �p�   �_�       ���  ����  Ɲ��  �> ���  L?    �A�  ����  ��O�  �? ���  �Z�  �? ���  ����  Ɲ��  �? ���  ���  �? ���  "@ �F�  ����  ��T�  s@ ���   � �_�  �@ ��  ��   V��  �@   �`�   �T�  �@ �`�   �_�           �l�  ,��  �� �z�  �@ ���  ,��  ����  �@ ��  ���  A ���  %A �F�  F�(�  ��T�  ]A �F�   � �_�  {A ��  O�   V��  �A   ���   �T�  �A ���   �_�        �Mz  ��   %2 �[z  �A �4z  ��   	��Bz  �A �z  ��   	-�$z  �A    ��  ־   E� ��  B ���  )B ���  ־   ���  B ���  =B   ��  �@�  F� ���  RB �4z  �   	#� �Bz  RB  ��}  �h�  	#��}  �B ��}  �B �3���  �Ruc   ���  ���  (- �Ȍ  �B ���  �B �!���   �Mz  S�   2� �[z  eC �4z  S�   	��Bz  eC �z  S�   	-�$z  eC    �l�  ��   �� �z�  zC ��  ��   �� ��   �����   ���  :���  �b ���  �C ��  D���  ��,�  �C �D�   : �7�  �{  M�   B�+{  �5{  �C   � �+   �,�  D � �+   �7�      ���  Z�   �� �ˆ  D ���  JD �g���   �l�  ��Ќ  �� �z�  �D ��  ��   �� ��   �����   ��  ��   FS ���  ud��4z  ��   	# �Bz  ud� ��}  ��   	#��}  �D ��}  �D �����  �Ruc   ��+E �6�j  ���3   ���Ge  �u  �w  �x  ]u  �B  � � �h  ��  ��|  ��?  ��h  ��?  �$  �� ��*  �� �__v ��  �u  �w  �x  �� G�  ��7   � W �� ��� ��� ��� ��� ��� � ����
  �@  ��|   �o  �h  ��  ��e  ��?  ���h  ��?  ��$  � ���*  �" ��__v �' � �� �&   ��� E �� E �� 3E �� �� �� RE �0��
   �u  �w  �x  ��E  p��  �M �) ]T  k  �h  ��  ���|  rD6  ���h  rD6  ��$  r�) ���*  s�) ��__v s�) � ��  �) Tߠ  wks  T��  x�=  �ϴ  yia  �Z�ȱ  z�) ��k  {� qE   � �ԥ  |�j  �E �__c }y?  zF ��m  ��$  �'�  �u  WG ���  ��j  �G � �  ��t  H ���  ��t  I �Qr  ��t  yI ���  ��j  J �R'  ��c  �J �p�  ��!  �\���  ��t  gK ���  ��t  �K ��  �� ZL � �ڪ  �� �L ��T  �� �L �9�  ��j  wM �S�  �m� �M �}�  |�   zW ���  |N  �(�  ���  �~ �>�  J�2�  �N  �3�  �� �  �� �[�  �N �O�  �O �����   �l�  ��8�  �� �z�  "P ��  ��   �� ��   �����   ���  �   �! ���  �P ���   ���  )�   �U �ˆ  �P ���  �P �6���   ���  l�   �� ���  Q �X�  l�   	��}�  �p�  qQ �f�  Q   �:�  ��P�  �4 �m�  �Q �`�  �Q �[�  �Q �Q�  R ���&   � �{�  AR  �p�  �Q�  �R �[�  �R �`�  �R �m�  �p�  �{�  �R    ���  ����  �� ���  "S ��  ����  ��,�  DS �؍  � �7�  �{  ����  B�+{  �5{  bS   � �   �,�  vS � �   �7�      ���  ��  ��! �ˆ  �S ���  �S ���  ��  ԝ�  �S ��  �S �A�  �0�  �! �O�  �S �0�  �Z�  �S ���  �`�  ��  ���  �S �`�  ���  �S ���  �S �F�  ���  ��T�  @T ���  �  �_�  ^T ��  �   V��  �T   �0�   �T�  �T �0�   �_�       ���  '���  Ɲ��  �T ���  :U    �A�  �Ȏ  ��O�  �U �Ȏ  �Z�  �U ���  �Ȏ  Ɲ��  �U �Ȏ  ���  �U ���  0V �F�  �� �  ��T�  uV ���   �! �_�  �V ��  ��   V��  �V   �p�   �T�  �V �p�   �_�           �l�  ��   5" �z�  �V ��  ��   �*" ��   �����   ��  �" �__q 
m� �I  ��   �m  W �`  8W �S  XW ���Bg   ���  ��   ��" �Ȍ  zW ���  �W �����   ���   �0�  O# ���  �W ��  
�X�  ��,�   X �x�  '# �7�  �{  ���  B�+{  �5{  X   ���   �,�  2X ���   �7�      ���  #���  w% �ˆ  EX ���  gX ���  #���  ԝ�  EX ��  gX �A�  #�Џ  ��$ �O�  gX �Џ  �Z�  �X ���  #� �  �v$ ���  gX � �  ���  �X ���  �X �F�  #� �  ��T�  �X �8�  M$ �_�  Y ��  ,�   V��  DY   � �   �T�  WY � �   �_�       ���  =�P�  Ɲ��  jY ���  �Y    �A�  /�h�  ��O�  4Z �h�  �Z�  VZ ���  /�h�  Ɲ��  4Z �h�  ���  VZ ���  �Z �F�  ����  ��T�  �Z ���   J% �_�  [ ��  ��   V��  +[   ���   �T�  >[ ���   �_�           �l�  ����  �C& �z�  Q[ ���  ����  ����  Q[ ���  ���  s[ ���  �[ �F�  ��А  ��T�  �[ ���   & �_�  �[ ��  ��   V��  	\   �`�   �T�  \ �`�   �_�        �Mz  C�   %�& �[z  /\ �4z  C�   	��Bz  /\ �z  C�   	-�$z  /\    ��  v�   E�& ��  �\ ���  �\ ���  v�   ���  �\ ���  �\   ��  ���  Fb' ���  �\ �4z  ��   	#)' �Bz  �\  ��}  ���  	#��}  �\ ��}  :] �����  �Ruc   ���  ��0�  (�' �Ȍ  X] ���  l] �����   �Mz  ��   2�' �[z  �] �4z  ��   	��Bz  �] �z  ��   	-�$z  �]    �l�  0�   �3( �z�  �] ��  <�   �(( ��   �<���   ���  ��H�  ��( ���  ^ ��  ��`�  ��,�  F^ ���   �( �7�  �{  ��   B�+{  �5{  d^   ���+   �,�  x^ ���+   �7�      ���  ��   ��( �ˆ  �^ ���  �^ �����   �l�  P�x�  �D) �z�  _ ��  c�   �9) ��   �\���   ��  �   F�) ���  ud��4z  �   	#�) �Bz  ud� ��}  �   	#��}  ;_ ��}  h_ �%���  �Ruc   ���+E ���j  ��3   �.�Ge  �u  �w  �x  ]u  /C  * T* �h  ��  ��|  ��?  ��h  ��?  �$  �T* ��*  �Y* �__v �^*  �u  �w  �x  ��) �  0�7   �* �* �* ��* ��* ��,* ��9* ��F* � �^�,  �W@  p�|   ��* �+ �h  ��  ��e  ��?  ���h  ��?  ��$  ��+ ���*  ��+ ��__v ��+ � ��) ��&   ��F* {_ �9* �_ �,* �_ �* �* �* �_ ���,   �u  �w  �x  �*F  ���  ��+ O: ]T  7   �h  ��  ���|  rD6  ���h  rD6  ��$  rO: ���*  sT: ��__v sY: � ���  D: Tߠ  w�s  T��  x�=  �ϴ  yia  �Z�ȱ  z^: ��k  {c, �_ i, ), �ԥ  |�j  T` �__c }y?  �` ��m  ��$  �'�  �u  �a ���  ��j  /b � �  ��t  sb ���  ��t  �c �Qr  ��t  �c ���  ��j  ud �R'  ��c  ne �p�  ��!  �\���  ��t  �e ���  ��t  ;f ��  �W- �f , �ڪ  �W- g ��T  �, ng �9�  ��j  �g �S�  �m� h �}�  ��   z�- ���  �h  �(�  	���  ��- �>�  J�2�  -i  �3�  4�ȑ  �. �[�  Li �O�  j �D���   �l�  R���  �`. �z�  �j ��  d�   �U. ��   �^���   ���  ��   ��. ���  �j ����   ���  ��   ��. �ˆ  k ���  6k �����   ���  ��   �
/ ���  pk �X�  ��   	��}�  �p�  �k �f�  pk   �:�  ,���  ��/ �m�   l �`�   l �[�  Ll �Q�  �l �,�&   `/ �{�  �l  ��  �Q�   m �[�   m �`�  Hm �m�  ��  �{�  hm    ���  a�8�  �10 ���  �m ��  t�`�  ��,�  �m ���  	0 �7�  �{  }���  B�+{  �5{  �m   ���   �,�  �m ���   �7�      ���  ����  �Y2 �ˆ  �m ���  n ���  ����  ԝ�  �m ��  n �A�  ��ؒ  �1 �O�  n �ؒ  �Z�  <n ���  ���  �X1 ���  n ��  ���  <n ���  ^n �F�  ��(�  ��T�  �n �@�  /1 �_�  �n ��  ��   V��  �n   ���   �T�  
o ���   �_�       ���  ��X�  Ɲ��  o ���  �o    �A�  ��p�  ��O�  Ap �p�  �Z�  cp ���  ��p�  Ɲ��  Ap �p�  ���  cp ���  �p �F�  +���  ��T�  �p �+�   ,2 �_�  q ��  4�   V��  ,q   ���   �T�  ?q ���   �_�           �l�  �   �2 �z�  Rq ��  �   ��2 ��   ����   ���  �2 �__q 
m� �I  @�   �m  q �`  �q �S  �q �P�Bg   ���  +�   �$3 �Ȍ  �q ���   r �;���   ���  ��ؓ  �3 ���  Mr ��  �� �  ��,�  or � �  �3 �7�  �{  ��8�  B�+{  �5{  �r   �P�   �,�  �r �P�   �7�      ���  ��P�  �5 �ˆ  �r ���  �r ���  ��P�  ԝ�  �r ��  �r �A�  ��x�  �5 �O�  �r �x�  �Z�  �r ���  ����  ��4 ���  �r ���  ���  �r ���  s �F�  ��Ȕ  ��T�  ks ���  �4 �_�  �s ��  ��   V��  �s   ���   �T�  �s ���   �_�       ���  ����  Ɲ��  �s ���  +t    �A�  ���  ��O�  �t ��  �Z�  �t ���  ���  Ɲ��  �t ��  ���  �t ���  u �F�  �H�  ��T�  Ru ��   �5 �_�  pu ��  �   V��  �u   �`�   �T�  �u �`�   �_�           �l�  D�`�  ��6 �z�  �u ���  D�`�  ����  �u �`�  ���  �u ���  v �F�  ^�x�  ��T�  <v �^�   �6 �_�  Zv ��  c�   V��  xv   ���   �T�  �v ���   �_�        �Mz  ��   %7 �[z  �v �4z  ��   	��Bz  �v �z  ��   	-�$z  �v    ��  ��   ES7 ��  �v ���  w ���  ��   ���  �v ���  w   ��  ���  F�7 ���  1w �4z  �   	#�7 �Bz  1w  ��}  ���  	#��}  mw ��}  �w �3���  �Ruc   ���  0�ؕ  (�7 �Ȍ  �w ���  �w �A���   �Mz  s�   2W8 �[z  Dx �4z  s�   	��Bz  Dx �z  s�   	-�$z  Dx    �l�  ��   ��8 �z�  Yx ��  ��   ��8 ��   �����   ���  :��  �49 ���  �x ��  D��  ��,�  �x �D�   9 �7�  �{  M�   B�+{  �5{  �x   � �+   �,�  �x � �+   �7�      ���  Z�   �h9 �ˆ  �x ���  )y �g���   �l�  �� �  ��9 �z�  py ��  ��   ��9 ��   �����   ��  ��   F%: ���  ud��4z  ��   	#�9 �Bz  ud� ��}  ��   	#��}  �y ��}  �y �����  �Ruc   �	�+E �V�j  ���3   ���Ge  �u  �w  �x  ]u  oC  q: �: �h  ��  ��|  ��?  ��h  ��?  �$  ��: ��*  ��: �__v ��:  �u  �w  �x  �c: ��  ��7   ��: ); �q: ��{: ���: ���: ���: ���: � ����+  ��D  ��l   �A; y< �h  ��  ���|  ��?  �y ��h  ��?  ��$  �y< ���*  �~< ��__v ��< � �8�  T�P  ��#  �-  ��; �; T��  ��r  �v|  ��; �l�(�  �   �< �>�  ��2�  z  ��  �   �.< �4�  �(�  0z  �=�  ?�   �m< �K�  wz �U�  �z �?�   �c�  �z   �7��+   �u  �w  �x  ��@  `�|   ��< N= �h  ��  ��e  ��?  ���h  ��?  ��$  �N= ���*  �S= ��__v �X= � �c: }�&   ���: �z ��: �z ��: �z ��: �{: �q: { ����+   �u  �w  �x  �kF  ���	  �~= L ]T  0k  �h  ��  ���|  rD6  ���h  rD6  ��$  rL ���*  sL ��__v sL � �P�  L Tߠ  w�l  T��  x�=  �ϴ  yia  �Z�ȱ  z"L ��k  {+> 2{ 1> �= �ԥ  |�j  �{ �__c }y?  �{ ��m  ��$  �'�  �u  �| ���  ��j  m} � �  ��t  �} ���  ��t    �Qr  ��t  � ���  ��j  .� �R'  ��c  8� �p�  ��!  �\���  ��t  X� ���  ��t  ԁ ��  �? y� �= �ڪ  �? �� ��T  ��= �� �9�  ��j  �� �S�  �m� 
� �}�  ��   z�? ���  ��  �(�  ��p�  ��? �>�  J�2�  �  �3�  &���  ��? �[�  � �O�  ӆ �6���   �l�  D���  �(@ �z�  L� ��  V�   �@ ��   �P���   ���  w�   �R@ ���  �� ����   ���  ��   ��@ �ˆ  ܇ ���  �� �����   ���  ��   ��@ ���  8� �X�  ��   	��}�  �p�  �� �f�  8�   ���  $A �__q 
m� �I  x�   �m  Ո �`  � �S  9� ���Bg   ���  ��   �XA �Ȍ  h� ���  �� ����   ���  &���  �A ���  ͉ ��  4��  ��,�  � �(�  �A �7�  �{  =�@�  B�+{  �5{  �   � �   �,�  !� � �   �7�      ���  M�X�  D �ˆ  4� ���  V� ���  M�X�  ԝ�  4� ��  V� �A�  M���  �:C �O�  V� ���  �Z�  x� ���  M���  �C ���  V� ���  ���  x� ���  �� �F�  M�З  ��T�  � ��  �B �_�  	� ��  V�   V��  3�   �P�   �T�  F� �P�   �_�       ���  g� �  Ɲ��  Y� ���  ��    �A�  Y��  ��O�  #� ��  �Z�  E� ���  Y��  Ɲ��  #� ��  ���  E� ���  t� �F�  ��P�  ��T�  �� ���   �C �_�  ׌ ��  ��   V��  �   ���   �T�  � ���   �_�           �l�  ��   YD �z�  '� ��  ��   �ND ��   �����   �:�  ��h�  ��D �m�  T� �`�  � �[�  �� �Q�  Í ���  �D �{�  �  ���  �Q�  ,� �[�  L� �`�  p� �m�  ���  �{�  ��    ���  ����  �|E ���  Ď ��  ���  ��,�  � ��  TE �7�  �{  ��(�  B�+{  �5{  �   �@�   �,�  � �@�   �7�      ���  ��@�  ��G �ˆ  +� ���  M� ���  ��@�  ԝ�  +� ��  M� �A�  ��h�  ��F �O�  M� �h�  �Z�  o� ���  ����  ƣF ���  M� ���  ���  o� ���  �� �F�  ����  ��T�  � �Й  zF �_�   � ��  ��   V��  *�   �p�   �T�  =� �p�   �_�       ���  ��  Ɲ��  P� ���  �    �A�  � �  ��O�  �� � �  �Z�  �� ���  � �  Ɲ��  �� � �  ���  �� ���  � �F�  �8�  ��T�  =� ��   wG �_�  [� ��  �   V��  ��   ��   �T�  �� ��   �_�           �l�  !�P�  �pH �z�  �� ���  !�P�  ����  �� �P�  ���  ڒ ���  	� �F�  s�p�  ��T�  N� �s�   FH �_�  l� ��  |�   V��  ��   ���   �T�  �� ���   �_�        �Mz  ��   %�H �[z  �� �4z  ��   	��Bz  �� �z  ��   	-�$z  ��    ��  ��   EI ��  � ���  '� ���  ��   ���  � ���  ;�   ��  ����  F�I ���  P� �4z  ��   	#VI �Bz  P�  ��}  ����  	#��}  �� ��}  Ȕ �i���  �Ruc   ���   �К  (�I �Ȍ  � ���  �� ����   �Mz  @�   2J �[z  @� �4z  @�   	��Bz  @� �z  @�   	-�$z  @�    �l�  �   �`J �z�  U� ��  �   �UJ ��   ����   ���  ���  ��J ���  �� ��  �� �  ��,�  �� ���   �J �7�  �{  ��   B�+{  �5{  ܕ   �P�   �,�  � �P�   �7�      ���  ��   �,K �ˆ  � ���  2� �����   �l�  ��  �qK �z�  y� ��  #�   �fK ��   ����   ��  ��   F�K ���  ud��4z  ��   	#�K �Bz  ud� ��}  ��   	#��}  �� ��}  �� �����  �Ruc   ���+E �#�j  ���3   ���Ge  �u  �w  �x  ]u  �C  5L �L �h  ��  ��|  ��?  ��h  ��?  �$  ��L ��*  ��L �__v ��L  �u  �w  �x  �'L ��  ��7   ��L �L �5L ��?L ��LL ��YL ��fL ��sL � ��]=  ��@   �|   �M �M �h  ��  ��e  ��?  ���h  ��?  ��$  ��M ���*  ��M ��__v ��M � �'L =�&   ��sL � �fL � �YL � �LL �?L �5L :� �`�]=   �u  �w  �x  ��F  ���	  ��M |\ ]T  )k  �h  ��  ���|  rD6  ���h  rD6  ��$  r|\ ���*  s�\ ��__v s�\ � �0�  q\ Tߠ  w�s  T��  x�=  �ϴ  yia  �Z�ȱ  z�\ ��k  {�N Y� �N VN �ԥ  |�j  �� �__c }y?  � ��m  ��$  �'�  �u  �� ���  ��j  R� � �  ��t  �� ���  ��t  �� �Qr  ��t  � ���  ��j  �� �R'  ��c  �� �p�  ��!  �\���  ��t  Ԝ ���  ��t  9� ��  ��O ѝ JN �ڪ  ��O )� ��T  �JN �� �9�  ��j  � �S�  �m� s� �}�  ��   z�O ���  *�  �(�  ��X�  �P �>�  J�2�  l�  �3�  ��x�  �HP �[�  �� �O�  L� �����   �l�  ����  ��P �z�  Ţ ��  �   ��P ��   ����   ���  <�   ��P ���  &� �L��   ���  V�   ��P �ˆ  H� ���  j� �c���   ���  ��   �7Q ���  �� �X�  ��   	��}�  �p�  � �f�  ��   �:�  ����  ��Q �m�  4� �`�  T� �[�  �� �Q�  �� ���&   �Q �{�  �  ���  �Q�  A� �[�  U� �`�  m� �m�  ���  �{�  ��    ���  9�؛  �^R ���  �� ��  K��  ��,�  �� �(�  6R �7�  �{  T�@�  B�+{  �5{  ԥ   ���   �,�  � ���   �7�      ���  d�X�  ��T �ˆ  �� ���  � ���  d�X�  ԝ�  �� ��  � �A�  d���  ��S �O�  � ���  �Z�  ?� ���  d���  ƅS ���  � ���  ���  ?� ���  a� �F�  d�М  ��T�  �� ��  \S �_�  Ц ��  m�   V��  ��   ���   �T�  � ���   �_�       ���  ~� �  Ɲ��   � ���  ��    �A�  p��  ��O�  D� ��  �Z�  f� ���  p��  Ɲ��  D� ��  ���  f� ���  �� �F�  [�P�  ��T�  � �[�   YT �_�  � ��  d�   V��  /�   ���   �T�  B� ���   �_�           �h�  �T �__q 
m� �I  ��   �m  U� �`  }� �S  �� ���Bg   ���  ��   �U �Ȍ  �� ���  �� �����   ���  S���  �U ���  $� ��  a���  ��,�  F� �Н  xU �7�  �{  j��  B�+{  �5{  d�   ���   �,�  x� ���   �7�      ���  z� �  �W �ˆ  �� ���  �� ���  z� �  ԝ�  �� ��  �� �A�  z�(�  ��V �O�  �� �(�  �Z�  Ϫ ���  z�X�  ��V ���  �� �X�  ���  Ϫ ���  � �F�  z�x�  ��T�  B� ���  �V �_�  `� ��  ��   V��  ��   � �   �T�  �� � �   �_�       ���  ����  Ɲ��  �� ���  �    �A�  ����  ��O�  j� ���  �Z�  �� ���  ����  Ɲ��  j� ���  ���  �� ���  �� �F�  ����  ��T�  � ���   �W �_�  *� ��  ��   V��  T�   �0�   �T�  g� �0�   �_�           �l�  ��   X �z�  z� ��  ��   �X ��   �����   �l�  t��  ��X �z�  �� ���  t��  ����  �� ��  ���  ɭ ���  � �F�  ��(�  ��T�  #� ���   �X �_�  A� ��  ��   V��  _�   ��   �T�  r� ��   �_�        �Mz  ��   %1Y �[z  �� �4z  ��   	��Bz  �� �z  ��   	-�$z  ��    ��  ��   E�Y ��  ۮ ���  � ���  ��   ���  ۮ ���  �   ��  ��@�  F�Y ���  � �4z  ��   	#�Y �Bz  �  ��}  ��h�  	#��}  T� ��}  �� �����  �Ruc   ���  ���  (,Z �Ȍ  �� ���  ï �!���   �Mz  P�   2�Z �[z  � �4z  P�   	��Bz  � �z  P�   	-�$z  �    �l�  ��   ��Z �z�  � ��  ��   ��Z ��   �����   ���  ���  �a[ ���  2� ��  ���  ��,�  a� ��   9[ �7�  �{  �   B�+{  �5{  �   ���   �,�  �� ���   �7�      ���  ,�   ��[ �ˆ  �� ���  հ �9���   �l�  ��П  ��[ �z�  � ��  ��   ��[ ��   �����   ��  .�   FR\ ���  ud��4z  .�   	#\ �Bz  ud� ��}  4�   	#��}  V� ��}  �� �C���  �Ruc   ���+E �3�j  �n�3   �L�Ge  �u  �w  �x  ]u  �C  �\ �\ �h  ��  ��|  ��?  ��h  ��?  �$  ��\ ��*  ��\ �__v ��\  �u  �w  �x  ��\ %�  P�7   �] V] ��\ ���\ ���\ ���\ ���\ ���\ � �~��M  ��@  ��|   �n] ^ �h  ��  ��e  ��?  ���h  ��?  ��$  �^ ���*  �!^ ��__v �&^ � ��\ ��&   ���\ �� ��\ �� ��\ �� ��\ ��\ ��\ ݱ ����M   �u  �w  �x  �ڥ  ���   �a^ �1�  ���   B�<�  �I�  ��  �U  $=n^  7k  ��   $>n^ �B  $?n^ ��  $E�^  Bk  �B   $F�^ �C  $G�^ �e  $H�^ �8  $I�^ ��  $J�^ �

  $X�^  Mk  ��  $Y�^ ��
  $Z�^ ��   $`_ Xk  ��  $f+_  ck  ��  $g+_ ��  $h+_ ��  $nW_  nk  ��	  $oW_ ��  $pW_ �H  $v�_  yk  �`  $w�_ �w  $x�_ �   $y�_ �~  $�_  �k  �   $��_ ��  $��_ �  $��_ ��   $��_ ��  $��_ ��	  $��_ ��  $�`  �k  �  $�` �  $�` ��  $�` ��  $�U`  �k  ��  $�U` ��  $�U` ��  $�U` �m  $��`  �k  �	  $��` �2	  $��` ��  $��` �9  $��` �[  $��`  �k  �J  $��` ��  $��` �7  $��` ��  $�a  �k  �I	  $�a �$	  $�a ��   $�9a  �k  �N  $�9a �p  $�Xa  �k  ��  $�Xa �:  $�Xa ��  $�Xa �d   $�Xa ��  $ɞa  �k  �  $ʞa ��  $˞a ��	  $��a  �k  ��  $��a �  $��a  �k  ��  $��a ��  $��a ��  $��a �+  $�"b  �k  ��  $�"b ��   $�"b �  $�Nb  l  ��
  $�Nb ��  $�Nb �  $�zb  l  �   $�zb �F  $�zb ��  $�b  l  ��  $��b ��  $��b �D  %O�b  2l  ��  %P�b �1  %Q�b ��  %W�b  =l  �^  %X�b ��  &3c  Hl  ��  &4c ��   &8<c  Sl  ��  &9<c �l	  &=[c ^l  �N  &>[c �^  &?[c �L  &@[c �a  &D�c il  �B  &E�c ��	  &F�c �  &G�c �  &H�c �y  &I�c ��  ' �c  tl  ��  '!�c �j\  �u  �E�d;  H�  �E�m?  ��  �E�G  l�  �E��M  T�  �E�.  ��  B	�,.  +�  �E��(  �  C	��(  ��  �E�:Y  ��  �E�@3  �  A	��3  �  @	�64  3�  �E��7  ��  �E��R  ��  �E�lT  �  �E�e  0�Ӫ  e 0l   �  0�1  #e 0l   ��d  0l  Ae 0l  l  )l   v�-  �>  Y  [e 0l   �O2  Y2  7   se �j   0�  0��  0l  �e �   ��  ��  0l  �e 0l   ��  ��  �  �j  �e k  �j  �j   f�q  1h�j  �e �j   f�e  1r�j  �e �j   f܉  1+�j  f �j   fb  1^�j  "f �j   f��  1��j  7f �j   fWe  1|�j  Lf �j   f�d  1��j  af �j   f�e  1J�j  vf �j   f�  15�j  �f �j   f��  1��j  �f �j   �mw  ww  �j  �f �j  �j   ���  0l  �f l  �f �f %    �f q  2 �f �f �  ���  0l  0�  0��  0l   g �   �us  s  0l  Bg 0l  �j  7    ��`  �`  0l  l  �j  7     �   �5  ��  Y�  �V  ��      �  std  ,  %  0G�  c_� ��  �?  ��  K  \�   L   ��  qx   ~   	$   ��  s�   �   	$  
*   W  y�   	$  	�    U   >�  \  �   ��  q�   �   	f   ��  s�   �   	f  
l   W  y  	f  	�    �   %�  e �  &  7    $   Ey  �  $,?   -J   K  :�  �e  =?   � ?�  "  @�  �4  A  �J  B  �A  O�  �  	   �A  Q�  �  	  
   �A  V�  �  	  	�   �
 Y51  d  �    	  
|   �
 ]�R  p    &  	  
�   � c?  d  >  N  	  
X  
�   _ m.   b  r  	  
d  
X   �3  q89  X  �  �  	   .E  ��3  �  �  	  
d  
   �(  ��(  �  �  	  
d   _Tp �   L  :�  :s  �e  =?   � ?0  "  @=  �4  AH  �J  BN  �A  O:  @  	T   �A  QP  [  	T  
Z   �A  Vk  v  	T  	�   �
 YQ�  �  �  �  	`  
   �
 ]��    �  �  	`  
   � c��  �  �  �  	T  
�  
�   _ mQ�  �    	T  
�  
�   �3  q-�  �     &  	`   .E  ��  :  J  	T  
�  
N   �(  ���  ^  i  	T  
�   _Tp 6   �   �  o  �  �  �  �  �	  int (  #  �� �� �� 2*  7�  80    �  �  �    �  �    L  �  �  U   �   6    C  6  6  C  �  s  s  �     �  �  �  �  �  h  �     �  �  �  h  �  #  y   �  �  �  h  �  
�     *  �  �  h  �   T  [  	    h  �  #  y   @  *  9  h  �  
9   Z  h   L  V  h  V   $  >  �  �   �v    L  �  ~   �  �  h  V  __a s�   *    ��   �   ��  �  �  � �  � �   �  �  h  V  #  y   �  -�  0�   �    �  �  �   &  0  h  0   f    ��  @�   �P  Y  &  �  �   g  |  h  0  __a s|   l  Y  ��  P�   ��  �  g  � p  � �   �  �  h  0  #  y   �  �  `�   ��  �  �   �=   �7  ��  j�  �V  p�      g�  (  _� �7   �  �  8k  �{  k   ]�  k  \�   k  �D  !k  �3  "k  U>  #k  &�  $k  �  %k  �*  &k   ڡ  'q  $�U  (q  %TL  )q  &�I  *q  'Q  +q  (�C  ,q  )�J  -q  *1  .k  ,o(  /q  0�U  0q  1PL  1q  2�I  2q  3Q  3q  4�C  4q  5�J  5q  6 q  �  std % N'  5>   6N'  7z'  @4)  	%  0�=  �n  �b  �q  Fe  �h'  
�3  �=  �  G-  M-   �  eq �<-  S-    M-  M-   lt ��1  S-  !  M-  M-   ��  eF  h'  E  Z-  Z-  n   �K  �9  n  _  Z-   �(  
!  Z-  �  Z-  n  M-   1  �A  `-  �  `-  Z-  n   �5  �'  `-  �  `-  Z-  n   �3  �A  `-  �  `-  n  �   +  :  �  	  f-   �  �C   �P  �  (  M-   �B  $6  S-  G  f-  f-   eof (�:  �  ?  ,N0  �  f-    _� �7   �?  �%   K  	\  _)   �e  	_n  �4  	cl-  �J  	dr-  ��  	q�  �  �-   ��  	s�  �  �-  �-   W  	y�  �-  h'    �  �J  
pz  �B  
R  �   %  
k   �B  
A  �-  k  �-    �e  
y�  [V  
k  R  �G  
!   <  
x�  �4  
{�  �J  
|�  �J  
�*  `S  
�-  ~J  
�z  �J  
�  �%  
�  �K  
�R   I  
�R  :!  
��-   %H  
��  �   �3  2k  �G  7u'  t3  B�-  �'  
��O  �-  V  
��N  S-  [  a  �-   3  
�o+  S-  x  ~  �-   �P  
��O  �  �  �-   �M  
��P  �  �  �-   �,  
�-  �  �  �-  R   �+  
��R  k  �  �  �-   3  
�   k      �-  �-  �-   �/  !�B  �-  6  R  R  �-   �O  
�|6  I  T  �-  �-    (  ��6  h  s  �-  �-   !�   
�-  k  �  �  �-   "�1  o�*  k  �  �-  �-  R    !�A  
$n%  k  �  �  �-   !�A  
(�I  k  �  �  �-  k   !"A  
,�%  �-      �-   !�1  
2E)  �  -  3  �-   !�/  
6;&  �  K  Q  �-    �>  
:�>  e  k  �-   !S  
A:2  R  �  �  �-  R  o'    �#  
K�(  �  �  �-  R  R  o'   !9  
S>$  R  �  �  �-  R  R   !-U  
[�7  S-  �    �-  o'   #�5  
d�-  '  k  o'  R   #	1  
m�P  G  k  o'  R   #�3  
v\-  g  k  R  q   #nU  
��-  �  k  �  �   #nU  
�nG  �  k  �  �   #nU  
��   �  k  k  k   #nU  
�IP  �  k  o'  o'   �J  
�rR  h'  	  R  R    �=  ��H  	  /	  �-  R  R  R    V  �)  C	  I	  �-   $�'  
�D*  �-  %�0  
�j	  p	  �-   &�0  ��	  �	  �-  �-   �0  ��	  �	  �-  �-   �0  ��	  �	  �-  �-  R  R   �0  ��	  �	  �-  �-  R  R  �-   �0  �
  
  �-  o'  R  �-   �0  �*
  :
  �-  o'  �-   �0  �J
  _
  �-  R  q  �-   %�0  
"p
  {
  �-  h'   '�  
*,Q  �-  �
  �
  �-  �-   '�  
2�G  �-  �
  �
  �-  o'   '�  
=�%  �-  �
  �
  �-  q   'S� 
f�&  �       �-   'S� 
q�>  �    %  �-   (end 
y<  �  >  D  �-   (end 
�6;  �  ]  c  �-   'I 
��$  �  |  �  �-   'I 
��7  �  �  �  �-   '��  
�lC  �  �  �  �-   '��  
�CM  �  �  �  �-   'r 
��R  R  �  �  �-   '�K  
�r5  R      �-   '�3  
�j=  R  6  <  �-   )�� �  Q  a  �-  R  q   )�� 
��F  v  �  �-  R   'I  
v  R  �  �  �-   )�E  �|U  �  �  �-  R   )�1  
-�  �  �  �-   '�� 
5�?  S-  �  �  �-   '�:  
D�6  �      �-  R   '�:  
UW  �  7  B  �-  R   (at 
k
/  �  Z  e  �-  R   (at 
��7  �  }  �  �-  R   '�F  
��/  �-  �  �  �-  �-   '�F  
�k:  �-  �  �  �-  o'   '�F  
��H  �-  �  �  �-  q   '@  DA:  �-      �-  �-   '@  U�1  �-  1  F  �-  �-  R  R   '@  )�D  �-  _  o  �-  o'  R   '@  
��*  �-  �  �  �-  o'   '@  �6  �-  �  �  �-  R  q   )�G  
-aN  �  �  �-  q   *�3  �b*  �-  �  �  �-  �-   '�3  
^ 2  �-    -  �-  �-  R  R   '�3  �=  �-  F  V  �-  o'  R   '�3  
z�T  �-  o  z  �-  o'   '�3  
� @  �-  �  �  �-  R  q   )� 
��E  �  �  �-  �  R  q   '� 
�\+  �-  �  �  �-  R  �-   '� 
�u>  �-    )  �-  R  �-  R  R   '� g|=  �-  B  W  �-  R  o'  R   '� 
"�@  �-  p  �  �-  R  o'   '� 
9k<  �-  �  �  �-  R  R  q   '� 
K�'  �  �  �  �-  �  q   'bL  
d�R  �-  �     �-  R  R   'bL  
t�2  �    $  �-  �   'bL  �L&  �  =  M  �-  �  �   '�%  
�9F  �-  f  {  �-  R  R  �-   '�%  
�|<  �-  �  �  �-  R  R  �-  R  R   '�%  ��T  �-  �  �  �-  R  R  o'  R   '�%  
��A  �-  �    �-  R  R  o'   '�%  
b>  �-  -  G  �-  R  R  R  q   '�%  
3%  �-  `  u  �-  �  �  �-   '�%  
'V7  �-  �  �  �-  �  �  o'  R   '�%  
<�+  �-  �  �  �-  �  �  o'   '�%  
Q'S  �-  �  	  �-  �  �  R  q   '�%  
vj.  �-  "  <  �-  �  �  k  k   '�%  
��9  �-  U  o  �-  �  �  o'  o'   '�%  
�C  �-  �  �  �-  �  �  �  �   '�%  
�>/  �-  �  �  �-  �  �  �  �   !�?  ��&  �-  �    �-  R  R  R  q   !�1  �O  �-    9  �-  R  R  o'  R   ,)  
�z-  k  ]  R  q  �-   ++E  �3J  k  �  R  q  �-   '�5  ��)  R  �  �  �-  k  R  R   )n	 @D  �  �  �-  �-   'W�  
�6  o'  �  �  �-   '�A  
%�A  o'      �-   '��  
,Z5  }  %  +  �-   '�(  �;  R  D  Y  �-  o'  R  R   '�(  
I�%  R  r  �  �-  �-  R   '�(  
X�5  R  �  �  �-  o'  R   '�(  �^   R  �  �  �-  q  R   '�(  
v�S  R  �  �  �-  �-  R   '�(  	K  R    +  �-  o'  R  R   '�(  
�o?  R  D  T  �-  o'  R   '�(  J5  R  m  }  �-  q  R   'NW  
��Q  R  �  �  �-  �-  R   'NW  /�I  R  �  �  �-  o'  R  R   'NW  
��,  R  �  �  �-  o'  R   'NW  
��;  R    &  �-  q  R   '�S  
��I  R  ?  O  �-  �-  R   '�S  >T?  R  h  }  �-  o'  R  R   '�S  
05  R  �  �  �-  o'  R   '�S  
$S:  R  �  �  �-  q  R   '�>  
2hL  R  �  �  �-  �-  R   '�>  SUB  R    &  �-  o'  R  R   '�>  
Q�2  R  ?  O  �-  o'  R   '�>  _�K  R  h  x  �-  q  R   '�4  
qT  R  �  �  �-  �-  R   '�4  j�K  R  �  �  �-  o'  R  R   '�4  
��5  R  �  �  �-  o'  R   '�4  N.  R    !  �-  q  R   'U+  
�)  	  :  J  �-  R  R   '��  
�!1  h'  c  n  �-  �-   '��  ��T  h'  �  �  �-  R  R  �-   '��  ��O  h'  �  �  �-  R  R  �-  R  R   '��  �;.  h'  �  �  �-  o'   '��  ��B  h'    &  �-  R  R  o'   '��  ��,  h'  ?  Y  �-  R  R  o'  R     ,!T  q  -�E  �  -�F  �   .�&  .�7  	  �o  >-   �| Ch'  /Q  b�   �  /�F c�  /�R  d�  /3  e�  /�  f�  /�K  g�  /�@  h�   0all i�  ?1�� �d  :!  ��-   NF  �(.  �E  �n  p0  �(.  �%  �4.  2S  �:.  2�R  �:.  23  �:.  2�$  �:.  2�K  �:.  2�@  �:.  2�@  �E.   �4  �Z  �  �  �-    �=  y)  �  �  �-   3�� �    �-  [.  n   3��   %  �-  o'  n   3�� 5  @  �-  n   3N  P  [  �-  h'   3�� k  v  �-  [.    �  �U  �  �  �-  [.   !�&  �.  S-  �  �  �-    �F  &�;  �  �  �-  a.  �    �9  )�Q  �  �  �-  a.  P.    WR  ,`2      �-  a.  ".    �S  /=  3  C  �-  ".  ..   4e  7,  S  �-  ..  n    �$  �-   2OD  �-  2gP  �-  2�F  $�-  5< �  6�h  �ܧ  =    7id �C  �U  �n   2�I  ��-   �  �<?  �  �  .  .   8id �    .  .   9id �!  '  .   :4H  ��(  n  <  ".    �o  uS  Y  .   �o  ~i  t  .  
.   &�o  ��  �  .  o'   �o  ��  �  .  
.  o'  �   �o  ��  �  .  
.  
.  �   5  ��  �  .  h'   *�  ��*  
.      .  
.   *H�  ��N  2   /  5  .   *U  �9  S-  M  X  .  
.   *2  �t*  S-  p  {  .  
.   ;jP  �D  �  �  
.   <RD  �Q  
.  =�o  7�  �  .  �-   >�K  :�N  >�A  =�5  �K  @I  �  �  �    �,  CH<        .  
.  
.  �   �  �     �  � >	  �a  $�   rS  +�'  ?m�  ,`   I   ?��  -`   ?�4  .`   ?;�  /`   ?��  0`   ?� 1`    ?�� 2`   @@b  3`   @�e  4`    @�  5`    ?މ  6`   s�  'g.   <x.  =m.  >�.  @/  A/  B8/  CS/  Dn/  E�/  F�/  G�/  H�/  ד  �w!  ��  �y  � �k  �4  �l-  ,{�  k   v>0  wn0  {y0  ��0  ��0  ��0  ��0  �1  �21  �G1  �b1  �}1  ��1  ��1  ��1  ��1  ��1  �2  �32  �R2  Rg2  U�2  [�2  \�2  A�+   ��  8'  �   =    Bn�  �8'  B��  �S-  Bh�  ��   B��  ��   BF�  ��2  B>�  �q  B��  ��2  Cd�  ��2  C��  �q  Did -�  E��  �C'   F�b  �q  G�F ��"  #  �2  �2  S-  n   G�F �#  7#  �2  8'  �2  S-  n   His 1�c  S-  N#  ^#  �2  I   q   His p��  o'  u#  �#  �2  o'  o'  �2   *Oe  ��c  o'  �#  �#  �2  I   o'  o'   */�  �^�  o'  �#  �#  �2  I   o'  o'   'k�  ��  �"  �#  $  �2  �"   'k�  ,��  �2  !$  1$  �2  3  �2   �"  '��  <��  �"  O$  Z$  �2  �"   '��  M��  �2  s$  �$  �2  3  �2   '��  a�)  �"  �$  �$  �2  q   '��  |�  o'  �$  �$  �2  o'  o'  3   'g�  ��  q  �$  �$  �2  �"  q   'g�  ���  �2  %  1%  �2  �2  �2  q  k   'I�  �&�  �2  J%  P%  �2   <��  ���  �2  Ic�  5"  v%  �%  �2  h'   J�  ���  �"  "  �%  �%  �2  �"   J�  �_�  �2  "  �%  �%  �2  3  �2   J	�  }�  �"  "  �%  
&  �2  �"   J	�  ��  �2  "  +&  ;&  �2  3  �2   JKC  3�T  �"  "  \&  g&  �2  q   JKC  J��  o'  "  �&  �&  �2  o'  o'  3   J҉  d�  q  "  �&  �&  �2  �"  q   J҉  ~��  �2  	"  �&  	'  �2  �2  �2  q  k   ��  @�  '  "'  �2   K+3  W�3  1'  �2    W�  1�2  n  "   L)%  Kk  h'  h'  o'   Mint u'  q  NGT  P�'  >   �  �'  �  �  o  �	  �  qW  !h'    "�'  �  #  .  <�'  `  Dh'  �  W�'  �  _�'  �  eh'  t   mh'  a  uh'    ~h'  �  �h'  3  �h'  �  �h'  H  �h'  y  �h'    �h'  s  �h'  T   �h'  �  �h'  F  �h'  �  �h'  �  �h'    �h'  V  �h'  �  Os  N�'  �  V�'  \	  2h'  o  7h'  �  <h'  �  Ch'  �  h'  +)  PQpO qO !,)  R$   E-  	�  $,n  -y  K  :�*  �e  =n  � ?k  "  @o'  �4  Al-  �J  Br-  �A  O�)  �)  x-   �A  Q�)  �)  x-  ~-   �A  V�)  �)  x-  h'   *�
 Y51  w)  *  *  �-  �)   *�
 ]�R  �)  .*  9*  �-  �)   *� c?  w)  Q*  a*  x-  k)  %)   S_ m.   u*  �*  x-  w)  k)   *�3  q89  k)  �*  �*  �-   S.E  ��3  �*  �*  x-  w)  r-   S�(  ��(  �*  �*  x-  w)   T_Tp q   _)  UZD  �-  BF�  �k   F��  �L!  F�4  �b!  F� �W!  %��  �H+  N+  �/   G��  �_+  j+  �/  0   '*  ��}  +  �+  �+  0   'Ư  �?s  *+  �+  �+  0   '�F  �Ϭ  0  �+  �+  �/   '�F  ��  �*  �+  �+  �/  h'   'a�  �
�  0  ,  
,  �/   'a�   ��  �*  #,  .,  �/  h'   '�:  ,�  +  G,  R,  0  +   '�F  		n  0  k,  v,  �/  +   '(*  ��  �*  �,  �,  0  +   ' I  h�  0  �,  �,  �/  +   '�O  7k  �*  �,  �,  0  +   'WC  ]�  0  �,  -  0   ,{�  k  ,�  	   .8E  �*   �� �� �� R2*  7G-  V8�   W�  W�  �  �  �  W	  Wq  Wu'  _)  W�*  �*  �  W  �-    �    h'  h'    �  	    W  W�  W	  X7   �-  Y Y    �-  �-  o'  �  W-   -   �  W      ..  "   k  X".  E.  Y XP.  P.  Y V.  ".  W'   '   �-  �l  !%   j�  !#%   Ztm ,!,/  ,g  !.h'   �  !/h'  �  !0h'  ��  !1h'  ��  !2h'  ��  !3h'  ��  !4h'  �  !5h'  d�  !6h'   ��  !7%   $~�  !8o'  ( N\�  !>x.  Lѯ  !H&-  8/  m.  m.   L��  !Mm.  M/  M/   �.  L�  !Cm.  h/  h/   m.  L#�  !ak  �/  �/   �/  �.  L�� !fk  �/  �/   �/  m.  L��  !WM/  �/  �/   L[v  !\M/  �/  �/   L��  !R,   �/  k  ,   o'  �/   �*  W0  k  -  W�*  ["*  >0  �  "h'   \rem "h'   +  " 0  ["#@  n0  �  "$%    \rem "%%    A  "&I0  L� "�h'  �0  �0   �0  ]L�  ">&-  �0  o'   L�  "Hh'  �0  o'   L�  "I%   �0  o'   L�  "��(  �0  %)  %)  ,   ,   �0   1  ^h'  1  %)  %)   _div ">0  21  h'  h'   L    "�k  G1  o'   `�  " n0  b1  %   %    `�  ".h'  }1  o'  ,    `�  "\,   �1  �-  o'  ,    `3  ">h'  �1  �-  o'  ,    a�  "�1  �(  ,   ,   �0   Nk� "qh'  b�  "|�1  �'   L  "W&-  2  o'  4.   L  "f%   32  o'  4.  h'   L�  "g7   R2  o'  4.  h'   L?  "�h'  g2  o'   L��  #Eh'  �2  o'  o'   L��  #Uk  �2  h'   L��  #Ok  �2  k  o'   L��  #F,   �2  k  o'  ,    h'  `   Xq  �2  c�(  � "  H'  I   1$  �"  d  3  !3  eh  !3   .  f^�  G3  gw  �h'  g-�  �h'   d1%  U3  _3  eh  _3   �2  h;&  ��   �{3  �3  ih  _3  � j__c 3q  � h�&  ��   ��3  �3  ih  _3  � j__c d�"  �k�  dq  � da%   �3  �3  eh  �3  e#  �-   �2  l�3  Q�  p�W   �4  H4  m�3  � n���  n��=  o��p��n��.=   l�3  }�  ��   �c4  ~4  m�3  � n���3  q��B=   d�&  �4  �4  eh  _3  r�k  ~�2  r:�  ~�2  r�  q  r"y  k   l~4  ��  ��"   ��4  5  m�4  � m�4  �m�4  �m�4  �m�4  �n�W=   dg&  !5  O5  eh  _3  r�k  Jo'  r:�  Jo'  r"y  J3   l5  ��  ��"   �j5  �5  m!5  � m*5  �m65  �mB5  �n��W=   s	'   �   ��5  �6  th  _3  �� uب  vY�  C�2  ��}w �  �5  x__i Dn  �  y~4  d�0   F&6  z�4  ;� z�4  N� z�4  b� z�4  w� z�4  ��  w�  |6  {__c Oq  ��}|~4  ��   Pz�4  �� z�4  �� z�4  ǲ z�4  ݲ z�4  �   n��u=    s"'   ��   ��6  7  th  _3  � u8�  vY�  Z�2  ��}wX�  �6  x__i [n  #�  y5  ]�*   ]7  zB5  B� z65  U� z*5  j� z!5  }�  n��u=    }U  ='7   �'  }�   >'7  }B  ?'7  }�  EP7   �'  }B   FP7  }C  GP7  }e  HP7  }8  IP7  }�  JP7  }

  X�7   �'  }�  Y�7  }�
  Z�7  ~�   `�7  �'  }�  f�7   	(  }�  g�7  }�  h�7  }�  n 8   (  }�	  o 8  }�  p 8  }H  v)8   (  }`  w)8  }w  x)8  }   y)8  }~  ^8   *(  }   �^8  }�  �^8  }  �^8  }�   �^8  }�  �^8  }�	  �^8  }�  ��8   5(  }  ��8  }  ��8  }�  ��8  }�  ��8   @(  }�  ��8  }�  ��8  }�  ��8  }m  �!9   K(  }	  �!9  }2	  �!9  }�  �!9  }9  �!9  }[  �b9   V(  }J  �b9  }�  �b9  }7  �b9  }�  ��9   a(  }I	  ��9  }$	  ��9  }�   ��9   l(  }N  ��9  }p  ��9   w(  }�  ��9  }:  ��9  }�  ��9  }d   ��9  }�  �:   �(  }  �:  }�  �:  }�	  �G:   �(  }�  �G:  }  �d:   �(  }�  �d:  }�  �d:  }�  �d:  }+  �:   �(  }�  �:  }�   �:  }  ��:   �(  }�
  ��:  }�  ��:  }  ��:   �(  }   ��:  }F  ��:  }�  �;   �(  }�  �;  }�  �;  }D  O=;   �(  }�  P=;  }1  Q=;  }�  Wf;   �(  }^  Xf;  }�  3�;   �(  }�  4�;  }�   8�;   �(  }�  9�;  }l	  =�;  )  }N  >�;  }^  ?�;  }L  @�;  }a  D�;  )  }B  E�;  }�	  F�;  }  G�;  }  H�;  }y  I�;  }�   ?<   )  }�  !?<  T   O�  �	e   ��  �	q   %�  �	}   ��  �	�   ��  �	�   J�  �	�   �  �	�   ��  �	�   ��  �	�   -�  �	�   �  �	�"  >�  �E�"  ��  �	W8'  
�e  $�Ӫ  .=  �(   �>  Y  B=  �(   
�  $�1  W=  �(   ��d  �(  u=  �(  %)  �(   ���  ��  h'  %)  %)  7     b#   �?  [�  ��  �V  ث      �  (  _� 	�7   �  �  �  
P   �  �  o  �	  pW  
 w   �  qW  
!�   int   
"�   �    
#�   #  Fd ~   .  <~   `  D�   �  W~   �  _�   �  e�   t   m�   a  u�     ~�   �  ��   3  ��   �  ��   H  ��   y  ��     ��   s  ��   T   ȉ   �  Љ   F  ׉   �  ��   �  �     �   V  �   >   �  s  NE   �  VE   \	  2�   o  7�   �  <�   �  C�   �  �   E   	\  �   gX  �   X\  &3  X\  X,H  	$Z  .�    	\ /E   	� 1  	Z  2,   	K]  3E   	�_  4,   	\W  5,   	�Z  6,   	-_  8g   	VY  9�  $	`  :�  (	�Y  ;�  ,	7_  <�  0	BY  =   4	b\  >�  8	\  ?�  <	7Y  @�  @	 Z  A  D	SX  B  H	n4 Dl   L	`  Fa  P	*5 Ga  T 
  a  �  ,   a   3  H  
  �  �  ,   a   �  m  
�   �  a    �    �  
  �  a   �  
�   �  a   �  
a  �  �  �  a   �  >   �    a     pO qO !  std $ �  @  %  0�=  �  �b  �>   Fe  �   �3  �=    �  �   O  eq �<-  �  �  �  �   lt ��1  �  �  �  �   ��  eF  �   �  �  �     �K  �9    �  �   �(  
!  �     �    �   1  �A  �  D  �  �     �5  �'  �  h  �  �     �3  �A  �  �  �    O   +  :  O  �  �   Z  �C   �P  Z  �  �   �B  $6  �  �  �  �   eof (�:  Z  ?  ,N0  Z  �    _� �7   5�  6  77  �?  �%   W  3�  �4  �$  q-  c=  o'  �5   �%  � �8  �X)  ��%  ��  �aO  �Y=  � P  �� �C  ��wS  ��O  � �?  ��5  �� 
$ g�  )W  �   �U  �A  �8  �P   EH  �� �4  �+  O   �7  (  �Q  G  �� ��  �R  �R   �-  �1  lO  �� b4 �	  u�  �  �I  H  W�  �  u�  �  �  _   t�  �  _  �      �9  i�   �N  �+  !s0 B?  �  �  �  Q  �   "�P  �6  #d�  �c�  �    �   $�4  #  �  %dec #  $t-  #  %hex #  $r'  #  $< #   %oct #  @$� #  �&[)  #   &�%  "#   &�  &#   &dO  )#   &\=  ,#   &�P  /#    &�C  3#   @$zS  6#  �$�O  9#  J&�?  <#   �  J�  $�7  N9	  	  $(  Q9	  $�Q  V9	  $O  Y9	   %app lv	  �  %ate ov	  %in wv	  %out zv	  $�P  }v	   %beg ��	   �  %cur ��	  %end ��	   �8  I
  '�  T�	  
  �  �   �  �   "{'  E�
  (!T  >   )�E  C  *� �qP  e  B
  �    �Y  �
  '̾ ]b
  w
    �   �     "{'  E�
  (!T  >   )�E  C   �M  D  +Z  ��
  �
  �
  �  �    �B ��
  �
  �   ,��  �R�  �
     �  F  F  F   "�b  �>   ,��  +�  !  1  �  F  F   (!T  >   )�E  C   b(  ck  ev  f�  g�  h�  i�  j�  k�  l  m;  qU  rz  t�  u�  v�  x�  y  |  ~,  �>  �S  �m  �  ��  ��  ��  ��  �^  -(  -@�  �E  �  .tie -��  �  <  G  �  �   /`V    ]  h  �  �    aV  �y    �   (!T  >   )�E  C  0i3 ~P4  �  �  �  �   *3F  5u�  �  �  �  �    1�*  O6  �  6  6   1*  s�    �  �   ��  >  2�  ���  �  %  +  �   (!T  >   )�E  C     1	W  [�  ]  �  6   6  Ҿ �I
  3cin BT�  b  �  ��	  4��  C��  |  4M�  DH�  |  4A�  E<�  |   5$   ��  �  $,  -+  6U  AH  �  g  �    7��  I  g  �    W]  Z  8#`    !  ,  +  �    '$`  L<  G  +  �   (!T  >   )�E  C   69+  NH  t  g  �    7��  \�  g  �    9��  (!T  >   )�E  C    �� �� �� 52*  7�  -8<   :O  :  �    O  :�  �  8   	�{   �   	]�   �  	\�    �  	�D   !�  	�3   "�  	U>   #�  	&�   $�  	�   %�  	�*   &�   	ڡ   '>   $	�U   (>   %	TL   )>   &	�I   *>   '	Q   +>   (	�C   ,>   )	�J   ->   *	1   .�  ,	o(   />   0	�U   0>   1	PL   1>   2	�I   2>   3	Q   3>   4	�C   4>   5	�J   5>   6 1)%   K�  7  �   �   ;GT   PB  �  �  ! �     �   [  :�	  �^  "!  <Z  "1�  �   (  1aY  "��   �  �   =\  "C�   �  �   =xZ  "M�   �  �   1`  "��   �  �   =�^  "r�   �  �   =_X  "��     �     k  =�_  "��  ;  �  �   �   1�\  "��  U  �  �   =4Z  "�,   z  �  ,   ,   �   17`  "��  �  �  �  �   =>]  "	�   �  �  %   �    =�Z  "�   �  �  �   �  k  =�Y  " %   �  �   =�Y  "��     �   >\  "��   1�_  0�  ,  �   <�]  "W>  �   1D[  "T�   S  �   1�[  "a�   m  �  �   <�\  ")  �   ?Y@ "��  �  �   1�[  "   �  �  �  �   ,    ;�]  "i�  1D]  "w�  �  �   =}W  "��   �  �   �     5��  %g  -&�  4%�  )�    4��  *@�    4��  +�    4?�  -��  �  4��  .3�  �  4��  /��  �   H  @�  �  AXF  Ag  A\;  A�   BC�T  CH    @�  �  AXF  Ig  A\;  I�    �	    D#  �  �  Eh  �  Fl�  -�  BG'U  /�    �  �
  D�
    &  Eh  &  E#  Z   �    H  8A  T  Eh  T  E#  Z   +  DG  g  z  Eh  �  E#  Z   Dh  �  �  Eh  �   @�  �  I__c  �   �  D�
  �  �  Eh  &   J�  K�  #��  �    L__p #��   M�  #�  �  �   @�  %  L__a O6  L__b O6   @�  F  L__a s�  L__b s�      D�
  Z  �  Eh  &  F�  �F  F;�  �F  FP�  �F   D  �  �  Eh  &  FM�  +F  Fu�  +F   >  D  �  �  Eh  �   �  :]  :6  @C    L__a [  L__b [6   �  @Z  .  AXF  Ng  A\;  N�    D,  <  Q  Eh  T  L__f L�   R  D�  e  �  Eh  �  F�%  B�  BG'U  D�    Q  @t  �  AXF  \g  A\;  \�    H�  N�  �  Eh  �   _  �  
  D�	  �    Eh    E#  Z  E�!    A(  T�   �  �  I
  w
  DR
  3  Z  Eh  Z  E#  Z  E�!  _  A(  ]     �  N�  ���  ��  O�  ��  �P.  ����  U�  QE  �� R<  S�  ��P   MR�  T4�  P.  @�Щ  V�  QE  �� R<  U�  @��  MR�  T��  P.  ���  W7  QE  �� R<  U�  ��(�  MR�  T�  P�  �@�  [�  R  R�  Pz  �`�  Uv  Q�  ɳ T>� VY  -�!   U�  Qg  =� TF� W���   P%  ����  \  RN  R3  Pz  ����  ^�  Q�  Q� T�� VY  ��!   ^  Qg  }� T�� W��   P�  ���  ]x  R  R�  Pz  �Ȫ  UL  Q�  �� T*� VY  o�!   Un  Qg  � T�� W���   P�  ���  ^�  R  R�  Pz  ����  U�  Q�  �� T�� VY  N�!   U�  Qg  !� Tg� W ��   V�  �
   _  R�  R�  X�
   Y�    VW  �
   ``  Qn  5� Re  X�
   Y{  Z�  �
   EQ�  5� R�     V�  �
   c�  R�  R�  X�
   Y�    V�  !�   w�  Q�  K� R�  S�  !�   dQ�  K� R�    WN�:#  Wo�:#  W��:#  W��:#   [�  ��  ��%   �  r  O�  � P  ���  P^  \"  R  Um  ���  V\�  Rw  ]�  ^�  _�    _��d  `�  �   H�  { �  �  Eh  �  E#  Z   [r  C�  ��_   ��  0  Q�  r� P  ��(�    a"  R  Um  ��(�  Va�  Rw  ](�  ^�  ��    W �.
  W,�.
  W8�.
  WF�M#  bO�`#   c�  P�F  ��  d��  ��  � e@�  �  f�&  ��  �� ]`�  g]�  �[  �oP�  i�x�  ��  Q�  µ P  i���  P�  Q"  � R  Um  i���  VQ�  � Rw  ]��  ^�  �    hx�d  `�  uw  P1  ����  �-  RA  U  ����  8R  T��  V1  ��   �`  RA  S  ��   8R  T��  V1  ��   ��  RA  S  ��   8R  T��  T��T��T�W'��  W8��  WI��  WZ��  We��  W���    W��:#   iU  =�   �   i�   >�  iB  ?�  i�  E   �   iB   F  iC  G  ie  H  i8  I  i�  J  i

  Xf   �   i�  Yf  i�
  Zf  j�   `�  �   i�  f�   �   i�  g�  i�  h�  i�  n�   �   i�	  o�  i�  p�  iH  v�      i`  w�  iw  x�  i   y�  i~  '     i   �'  i�  �'  i  �'  i�   �'  i�  �'  i�	  �'  i�  ��     i  ��  i  ��  i�  ��  i�  ��   !  i�  ��  i�  ��  i�  ��  im  ��   ,  i	  ��  i2	  ��  i�  ��  i9  ��  i[  �+    7  iJ  �+   i�  �+   i7  �+   i�  �`    B  iI	  �`   i$	  �`   i�   ��    M  iN  ��   ip  ��    X  i�  ��   i:  ��   i�  ¦   id   æ   i�  ��    c  i  ��   i�  ��   i�	  �!   n  i�  �!  i  �-!   y  i�  �-!  i�  �-!  i�  �-!  i+  �b!   �  i�  �b!  i�   �b!  i  �!   �  i�
  �!  i�  �!  i  �!   �  i   �!  iF  �!  i�  ��!   �  i�  ��!  i�  ��!  iD  O"   �  i�  P"  i1  Q"  i�  W/"   �  i^  X/"  i�  3L"   �  i�  4L"  i�   8i"   �  i�  9i"  il	  =�"  �  iN  >�"  i^  ?�"  iL  @�"  ia  D�"  �  iB  E�"  i�	  F�"  i  G�"  i  H�"  iy  I�"  i�   #     i�  !#  kF�  "@�  k��  "B�  kz�  "D�  l>  Y  M#  �   m�  �  `#  �   n�   =N   F  � (�  �V  ��      �  std  �  ��  Y�$ _K   0     ��  c^   8     �  gq   K     %  0vj6  w�6  {�6  ��6  ��6  ��6  �7  �U7  �p7  ��7  ��7  ��7  ��7  �8  �)8  �48  �E8  �e8  ��8  ��8  G�  c_� �E4  �?  �h4  	K  	\~  
�   ��  	qE  K  �8   ��  	s[  f  �8  �8   W  	yr  �8  a4    "  
@�:  tr1 *�  ��  ��  Ic  ��   ��   `&    _1 h&  _2 i>  _3 jV  _4 kn  _5 l�  _6 m�  _7 n�  _8 o�  _9 p�  _10 q�  _11 r  _12 s.  _13 tF  _14 u^  _15 vv  _16 w�  _17 x�  _18 y�  _19 z�  _20 {�  _21 |  _22 }  _23 ~6  _24 N  _25 �f  _26 �~  _27 ��  _28 ��  _29 ��   g�   ��  X>  m�  a4   ��  XV  m�  a4   ]�  Xn  m�  a4   � X�  m�  a4   � X�  m�  a4   [ X�  m�  a4    X�  m�  a4   5 X�  m�  a4   ( X�  m�  a4  	 ( X  m�  a4  
 � X.  m�  a4   , XF  m�  a4   k X^  m�  a4   � Xv  m�  a4   y X�  m�  a4   N X�  m�  a4   3 X�  m�  a4   H X�  m�  a4   ` X�  m�  a4   � X  m�  a4   " X  m�  a4    X6  m�  a4    XN  m�  a4   � Xf  m�  a4   � X~  m�  a4   ��  X�  m�  a4   ��  X�  m�  a4   �  X�  m�  a4   ��  Xm�  a4    �  �  b	9  c�;  e<  f<  g3<  hI<  i_<  jt<  k�<  l�<  m�<  q�<  r
=  t)=  uI=  vo=  x�=  y�=  |�=  ~�=  ��=  ��=  ��=  �>  �%>  �I>  �T>  �i>  �=  �q  �b  �4  Fe  �a4  �3  �=  �  �>  �>   �  eq �<-  �8    �>  �>   lt ��1  �8  $  �>  �>   ��  eF  a4  H  �>  �>     �K  �9    b  �>   �(  
!  �>  �  �>    �>   1  �A  �>  �  �>  �>     �5  �'  �>  �  �>  �>     �3  �A  �>  �  �>    �   +  :  �    �>   �  �C   �P  �  +  �>   �B  $6  �8  J  �>  �>   eof (�:  �  ?  ,N0  �  �>    �:  Zo4  5�>  6�?  7�?  W  3 	   �4   �$   q-   c=   o'   �5    �%  �  �8  � X)  � �%  � �  � aO  � Y=  �  P  ��  �C  �� wS  � �O  �  �?  � �5  �� 
$ gY	   )W   �    �U   �A   �8   �P    EH  �� �4  ��	   O    �7   (   �Q   G  �� ��  ��	   �R    �-   �1   lO  �� !b4 �  "�9  i 	  "�N  ��	  #�P  ��  $�4  �	  �	  %dec �	  $t-  �	  %hex �	  $r'  �	  $< �	   %oct �	  @$� �	  �&[)  �	   &�%  "�	   &�  &�	   &dO  )�	   &\=  ,�	   &�P  /�	    &�C  3�	   @$zS  6�	  �$�O  9�	  J&�?  <�	  "�  JY	  $�7  N   �
  $(  Q   $�Q  V   $O  Y    %app l=  �	  %ate o=  %in w=  %out z=  $�P  }=   %beg ��   �	  %cur ��  %end ��   � H� �  �6   !�M  �  '�* �_e  �@  �  �  �@   #�b  ��4  (cb  �Pc      �@  a4   )Z  ��  '  2  �@  a4   (��  �R�  G  \  �@  �@  �@  �@   (��  +�  q  �  �@  �@  �@   *!T  �4  +�E  �   	�  5�  , 8�?   ,��  ;�8  � >�  �   @  @   -@�  Ad�   @  �      @  �6  �	  a4   -&�  Dx�   @    (   @  �?  �	   -&�  G(  @  @  P   @  a4  �	   -<_  JG�   @  h  n   @   -�  M��  �8  �  �  @   .fd P� a4  �  �   @   -QY  S� �?  �  �   @   � U�  �   @  a4   -�W  X" �  �  
   @  �6  �   -f [� �  "  <   @  �6  �  �6  �   -�W  _: �  T  d   @  �5  �   -09  b��  q  |  �   @  q  �	   -� e  a4  �  �   @   /��  h��  �  �   @    �^  -	9  � *�:  �  �>  b  !��  �  -�  ���  �8      �A   )�	 ��  '  2   B  a4   ( �< G  R   B  �   *!T  �4  +�E  �  -<_  ��  N  |  �   B   #��  S�  0Y /& �   B    �  1*  s 	  �   	   	   �  2%�  e �  �     3$   E04  �  $,  -  	K  :�  #�e  =  #� ?�5  #"  @�6  #�4  A�8  #�J  B�8  �A  OV  \  �8   �A  Ql  w  �8  �8   �A  V�  �  �8  a4   -�
 Y51    �  �  �8  .   -�
 ]�R  "  �  �  �8  :   -� c?    �     �8  
  47   4_ m.     $  �8    
   -�3  q89  
  <  B  �8   4.E  ��3  V  f  �8    �8   4�(  ��(  z  �  �8     5_Tp �4   �  D  3j�  E�  6� G \�    m�   \  E   J  K  ��  �^  7I�  �  8��  ��   9�  8B ��:  :��  �  )  ;  �   ;Q �� =  C  ;   <w �{�  �  W  ;    � ��  "   7� ��  8� �
;   7<  �"  =__C ��  =__L �Z  =__F �8  =__S �  >��  �A�  �  �  �  ;   >��  �j ;  �    ;   >��  �P ";       ;   �  :� �5  E  ;  
;  ";   :� �U  `  ;  ";   ��  �o
 �5  z     ?��  �5�  �  �5     � �q�  (;  �     ?\ �l�  �  (;     ��  ���  .;  �     ?q�  ���  �  .;     ��  ���  4;       ?d�  �� 4  4;     P�  �6�  :;  N     ?��  ���  i  :;     '�  �r�  @;  �  �  ;  F;   @� ��  �  ;  F;   *!T  �4  *�F  "   ��  F�  AF{2  AF�2  2   �  B M�  Bg N�8   8�  O04  8�	 P�5  8 �  R�:  7<  ]?2  :� bH  g  �;  �  a4  �8    H@   ,  ?M a�  �  �5    N@   ;"�  Sh �  �  �;   ;��  tm�  �  �  �;   ;D �9�  �  �  �;   ;. �j �  �  �;   ?� �� 
  �;   ?�  �h�     �;   ?� �s 6  �;   '�  �� T@  O  Z  �;  Z@   @� �k  v  �;  Z@   *!T  �4  *�F  "   >  �Z  �   89 ��;  8� ��;  7<  �?2  :
 ��  �  `@  �;  �;  f@   �  :	 �    `@  a4   '�  Q l@     +  `@  r@   @
 <  G  `@  r@   *!T  �4  *�F  "   ��  �8  �   8�A  ��5  7<  �?2  ��  �0�    �     :: ��  �  x@  �5    ~@   z  :9 ��  �  x@  a4   '�  �� �@  �  	  x@  �@   @: �  %  x@  �@   *!T  �4  *�F  "   �    �   8� �;  8"�  �8  7<  +?2  :��  -�  �  �@  �;    �8  �@   e  :��  >�  �  �@  a4   '�  G��  �@  �  �  �@  �@   @��  I�  �  �@  �@   *!T  �4  *�F  "   CW�  ^  D� �q/  A�}  A��  A�  
^   EY L;  F��  �l;  "�e  �  E[V  |
w  ]  "�J  �q/  "`S  �v/  "�4  �{/  "<  �  "� �  " �  "? Z  "��  8  "�    "~J  �  "�J  ,
�  G� q �8  &  �4   GE � �4  F  q;  ]   G��  (3�  �5  f  q;  ]   G��  ,| �8  �  w;  };       �  H� 4+ �  q;   H�  8s�  �  q;   G��  G� q;  �  q;       G! Jq�  q;    q;  �6     G3 O��  q;  2  q;  �6     Gm�  \)	 q;  R  q;  q;   (��  b��  g  |  �;      w;   G��  i   �     G�  mI�    �     Gx�  y�
 �;  �  �5    �;   GN �&�  �;  �  q;  q;  �;   G� �� �;  &  �;    �8  �;   G�  �u�  �;  P  �;      �;   G�  �w �;  u  �6    �;   G&�  � q;  �  q;  q;   G� �_ �;  �  �;  �6     G3�  �
�  �;  �  �;  �6     � ���    �  �6   :��  �	    �;  q;  �;   �  }�  �r�  �5  =  q;  �5   }�  ���  �5  f  q;      �5   ��  ���  �8  �  q;   ��  �� �8  �  q;   ��  �� �8  �  q;   ��  ���  q;  �  q;  q;   ��  �z�  q;  �  q;   ?(�  ��    q;  �;   ?S ���  #  q;  �;   ?��  I >  q;  a4   �J  ��  a4  ]  };  };   '�� 	�
 �8  v  |  �;   '��  � a4  �  �  �;  �;   @��  �  �  �;  �6  �;   @��  �  �  �;  �6    �;   @��  &�    �;  �6  �6  �;   @��  .  3  �;  �;  �;  �;   �  @��  4I  ^  �;  �;  �;  �;   |  @��  :t  �  �;  �4  �;   @��  L�  �  �;    �4  �;   @��  O�  �  �;  �;   @��  S�  �  �;  �;    �8  �;   @��  [      �;  �;  �;   @��  _#   .   �;  a4   '�  c&�  �;  G   R   �;  �;   (�1  m��  g   m   �;   (�G  t��  �   �   �;  �4   (H�  }��  �   �   �;   '�G  �� �4  �   �   �;   (��  ���  �   �   �;  �4   (� �V�  �   !  �;   '��  �B �4  !  !!  �;   (��  ���  6!  <!  �;   (�5  �_ Q!  \!  �;  �5   '�5  ���  ]  u!  �!  �;  ]  ]  �5   (��  �O�  �!  �!  �;   'W�  � �6  �!  �!  �;   '�
 ���  �6  �!  �!  �;   (P�  ��  �!  �!  �;   '�:  �:�  �4  "  ""  �;  ]   Iat ��  �4  :"  E"  �;  ]   'S� ��	 �  ^"  d"  �;   '��  �k �  }"  �"  �;   Iend  = �  �"  �"  �;   '��  � �  �"  �"  �;   'r � ]  �"  �"  �;   '�K  � ]  �"  �"  �;   '�3  � ]  #  #  �;   'I ��  �  7#  =#  �;   ' C
 �  V#  \#  �;   '��  #�	 �  u#  {#  �;   '� 'Q�  �  �#  �#  �;   '@  >/�  �;  �#  �#  �;  �6     '@  H� �;  �#  �#  �;  �6   '@  P� �;   $  $  �;  �6  �6   '@  Z+�  �;  )$  9$  �;  �  �   '@  go �;  R$  ]$  �;  �4   '@  q� �;  v$  |$  �;   '@  u��  �;  �$  �$  �;  �;   '@  ~T �;  �$  �$  �;    �4   (n	 �� �$  �$  �;  �;   G�%  �l	 q;  %  q;      q;   (� �D�  (%  8%  �;    �;   (� �R�  M%  b%  �;      �4   (� �� w%  �%  �;    �6     (� �� �%  �%  �;    �6   (� ���  �%  �%  �;    �4   (� �+�  �%  �%  �;     (� �N�  &   &  �;    �6  �6   (� ��  5&  J&  �;    �;  �;   (� ���  _&  t&  �;    �;  �;   (�%  � �&  �&  �;      �;   (�%  ��  �&  �&  �;      �6     (�%  �}�  �&  �&  �;      �4   (�%  	��  '  !'  �;      �6   (�%  	"�  6'  P'  �;      �6  �6   (�%  	��  e'  '  �;      �;  �;   (�%  	� �'  �'  �;      �;  �;   (�%  &	��  �'  �'  �;    �4   (�%  -	�  �'  �'  �;    �;   (�%  1	��  (  "(  �;    �6     (�%  5	��  7(  G(  �;    �6   (�%  9	��  \(  q(  �;    �6  �6   (�%  =	� �(  �(  �;    �;  �;   (�%  B	��  �(  �(  �;    �;  �;   (bL  H	e�  �(  �(  �;       (bL  R	 �(  
)  �;     '� W	� |  #)  3)  �;  �;  �;   '� ^	��  |  L)  a)  �;  �;    �4   '� d	��  |  z)  �)  �;  �;  �4   '� k	 |  �)  �)  �;  �;   '� r	� |  �)  �)  �;  �;  �6   '� y	}�  |  �)  *  �;  �;  �6     '� �	D |  *  3*  �;  �;  �6  �6   '� �	��  |  L*  a*  �;  �;  �;  �;   '� �	T |  z*  �*  �;  �;  �;  �;   (�%  �	��  �*  �*  �;  �;  �;  �;   (�%  �	  �*  �*  �;  �;  �;  �4   (�%  �	��  �*  +  �;  �;  �;  �6   (�%  �	� "+  <+  �;  �;  �;  �6     (�%  �	}�  Q+  k+  �;  �;  �;  �6  �6   (�%  �	��  �+  �+  �;  �;  �;  �;  �;   (�%  �	��  �+  �+  �;  �;  �;  �;  �;   (�%  �	%�  �+  �+  �;  �;  �;   (�%  �	��  ,  ,  �;  �;  �4   (�%  �	�  (,  8,  �;  �;  �6   (�%  �	(�  M,  b,  �;  �;  �6     (�%  �	��  w,  �,  �;  �;  �6  �6   (�%  �	��  �,  �,  �;  �;  �  �   (�%  �	 �,  �,  �;  �;  |  |   'bL  �	u |  �,  	-  �;  �;  �;   'bL  �	\�  |  "-  --  �;  �;   'U+  �	�   F-  V-  �;       'U+  �	G   o-  -  �;  |  |   'U+  �	�   �-  �-  �;  |   'U+   
f�    �-  �-  �;  �  �   'U+  

��    �-  �-  �;  �   '�(  
V�  ]  	.  .  �;  �4  ]   '�(  
� ]  2.  B.  �;  �6  ]   '��  %
� |  [.  a.  �;   '.�  )
z |  z.  �.  �;   'A /
��  �  �.  �.  �;   'x�  3
g�  �  �.  �.  �;   ' 7
��  �  �.  �.  �;  ]   Iend h
� �  �.  /  �;   'S� l
�  �  /   /  �;   '��  p
v �  9/  ?/  �;   'I t
�  �  X/  ^/  �;   *!T  �4  +�F  "   � ��  D
 ��0  8��  �   8F�  ��4  86�  ��8  7��  �  8� ��;  @��  ��/  �/  �;  �;     @��  ��/  0  �;  �;   @��  �0  +0  �;  �;    �4   'E � �4  D0  J0  �;   '�  �A�  �;  c0  n0  �;  �4   '*  �/ �0  �0  �0  �;   '�  �I�  �;  �0  �0  �;  �;   *!T  �4  *�F  "   � q�    !��  �0  *!T  �4   {/  C  F0   G^   C  7  :�  '1  J��  &�8  . K%1  L��  `2�  2  
�   #_� ;  � Aa1  g1  @   � w1  �1  @  a4  �	  E1   � ��1  �1  @  �?  �	  E1   )� {.1  �1  �1  @  a4   .fd m��  a4  �1  �1  @   -QY  w��  �?  2  2  @   *!T  �4  +�E  �   � $4  "   8o 8   7<  '"  =__C A�  =__L AZ  =__F A8  =__S A  >��  *��  ?2  �2  �2  @   >��  .��  @  �2  �2  $@   >��  2�  *@  �2  �2  @   ?2  :� 5�2  �2  $@    *@   ��  A��  �5  3     ?��  Al�  /3  �5     � A� 0@  I3     ?\ A� d3  0@     ��  A��  6@  ~3     ?q�  A� �3  6@     ��  AO�  <@  �3     ?d�  Aw�  �3  <@     P�  AE B@  �3     ?��  A��  4  B@     *!T  �4  *�F  "   2  �  �  Z  8   M�  Mo  M�  M�  M�  M�  M�	  Nint M(  M#  M�� M�� M�� 32*  7�4  K8q    M�  _�  �E4  �  !04  pW  ! >4  qW  !!a4    !"L4    !#o4  Os  "N�4  �  "V�4  PFd #�4  .  #<�4  `  #Da4  �  #W�4  �  #_�4  �  #ea4  t   #ma4  a  #ua4    #~a4  �  #�a4  3  #�a4  �  #�a4  H  #�a4  y  #�a4    #�a4  s  #�a4  T   #�a4  �  #�a4  F  #�a4  �  #�a4  �  #�a4    #�a4  V  #�a4  Q�4  M�  \	  $2a4  o  $7a4  �  $<a4  �  $Ca4  �  %a4  Q�4  R&*  j6  ,�  &a4   Srem &a4   +  & E6  R&#@  �6  ,�  &$h4   Srem &%h4   A  &&u6  1� &�a4  �6  �6   Q�6  T1�  &>}4  �6  �6   Q�6  �4  1�  &Ha4  �6  �6   1�  &Ih4  7  �6   1�  &��4  47  47  47  �4  �4  ;7   Q:7  UQA7  Va4  U7  47  47   Wdiv &j6  p7  a4  a4   1    &��5  �7  �6   X�  & �6  �7  h4  h4   X�  &.a4  �7  �6  �4   X�  &\�4  �7  �7  �6  �4   Q�7  M  X3  &>a4  8  �7  �6  �4   Y�  &)8  �4  �4  �4  ;7   Zk� &qa4  [�  &|E8  >4   1  &W}4  _8  �6  _8   Q�5  1  &fh4  �8  �6  _8  a4   1�  &gE4  �8  �6  _8  a4   1?  &�a4  �8  �6   \�4  \�6  Q�  \�  Q�  Q"  \~  �8  M�  a4  	\  '�4  gX  '�4  X\  (&9  X\  X(,):  ,$Z  (.�4   ,\ (/�4  ,� (1?6  ,Z  (2�4  ,K]  (3�4  ,�_  (4�4  ,\W  (5�4  ,�Z  (6�4  ,-_  (8H:   ,VY  (9g:  $,`  (:�:  (,�Y  (;�:  ,,7_  (<�:  0,BY  (=�:  4,b\  (>�:  8,\  (?�:  <,7Y  (@�:  @, Z  (A�:  D,SX  (B�:  H,n4 (D�4  L,`  (FB:  P,*5 (GB:  T V�8  B:  �4  �4  B:   Q9  Q):  V�8  g:  47  �4  B:   QN:  Va4  �:  B:  �8  a4   Qm:  V�8  �:  B:   Q�:  Va4  �:  B:   Q�:  VB:  �:  �6  �6  B:   Q�:  ]�:  B:   Q�:  ^)pO qO )!�:  ��  *!a4  Q�  Qq  Q  \�  Q^  \   Q�  Q�  Q�  Q�  \^  \  _�4  \;  `6    _E4  l;  `6  - \;  Q�  \�0  Q�  Q�0  Q�  \�  Q�  Q�  Q�0  Q�  Q�  Q  \  Qq;  \�0  \3  \^  \  Q�/  Q{/  \�0  Q�0  \{/  �^  +!�8  YZ  +1<  <   Q	9  1aY  +�a4  3<  <   X\  +Ca4  I<  <   XxZ  +Ma4  _<  <   1`  +�a4  t<  <   X�^  +ra4  �<  <   X_X  +�a4  �<  <  �<   Q�;  X�_  +��5  �<  �5  a4  <   1�\  +�<  �<  �6  �6   X4Z  +��4  
=  47  �4  �4  <   17`  +�<  )=  �6  �6  <   X>]  +	a4  I=  <  h4  a4   X�Z  +a4  d=  <  d=   Qj=  �;  X�Y  + h4  �=  <   X�Y  +�a4  �=  <   a\  +�a4  1�_  0�5  �=  �5   Y�]  +W�=  �6   1D[  +Ta4  �=  �6   1�[  +aa4  �=  �6  �6   Y�\  +)>  <   [Y@ +�%>  <  �5   1�[  +�a4  I>  <  �5  a4  �4   Z�]  +i<  1D]  +w�5  i>  �5   X}W  +�a4  �>  a4  <   \�  \�  Q�  Q�  \  �  8,�?  ,�{  ,�5   ,]�  ,�5  ,\�  , �5  ,�D  ,!�5  ,�3  ,"�5  ,U>  ,#�5  ,&�  ,$�5  ,�  ,%�5  ,�*  ,&�5   ,ڡ  ,'�4  $,�U  ,(�4  %,TL  ,)�4  &,�I  ,*�4  ',Q  ,+�4  (,�C  ,,�4  ),�J  ,-�4  *,1  ,.�5  ,,o(  ,/�4  0,�U  ,0�4  1,PL  ,1�4  2,�I  ,2�4  3,Q  ,3�4  4,�C  ,4�4  5,�J  ,5�4  6 1)%  ,K�5  �?  a4  �6   ZGT  ,P�?  Q�>  Q�  Q�  Q�  Q�  Q.1  Q4  \?2  Q2  \�2  QK2  QW2  Qc2  Qo2  \g  \,  \�  \4  Q�  \�  \�  \ 4  QZ  \�  \Z  \%4  Q8  \�  \8  \*4  Q�  Q�  b�  �@  �@  ch  �@   �@  Q�  b�  �@  �@  ch  �@  d__n �a4   �@  b  A  !A  ch  �@  c#  �8   e  8A  d__c  8A   �>  e+  `A  fhR  $`A  fmR  $eA   �>  �>  gJ  e�  �A  h__a s 	  h__b s 	   b2  �A  �A  ch  �@  f�  ��@  f;�  ��@  fP�  ��@   b\  �A  �A  ch  �@  fM�  +�@  fu�  +�@   Q�  b�  B  B  ch  B   �A  Q�  b  4B  GB  ch  GB  c#  �8    B  b�1   ZB  mB  ch  mB  c#  �8   @  iLB  n�  ��m   ��B  C  jZB  � k&B  �� �  |	C  l4B  "� k A  ���  ��B  lA  �� m�� n A  ��   ��B  lA  Ӷ o� p��d  o��o�� p�N   iLB   �   �.C  EC  jZB  � o�q+�.N   r&  &0�l   �D  s__r q;  �� s__i ]  4� t8�  u�  )�5  i� vX�  �C  w__l B�;  ��  vp�  �C  w__c 3�;  �� u�-  4q;  ˷ u��  5  �  xi�   w__f H�;  � y�T  I�4  �o   bQ1  D  'D  ch  mB   iD  Z�  ��   �BD  PD  jD  � o�� b2  ^D  �D  ch  GB  fQ  ��  z{�
 ��8  {8 ��8    bg1   �D  �D  ch  mB  |� �a4  |^F  ��	  |�a  �E1   i�D  _  ���   ��D  �E  j�D  � j�D  �j�D  �j�D  �nB  ��   �(E  lB  � p��n   kPD  "���  ��E  lgD  s� l^D  �� t��  }tD  �� ~�D  �A  0�   ��E  l�A  �� l�A  �� l�A  �  ��A  E�	   �l�A  6� l�A  6� l�A  6� l�A  ��    o��p��(  p"��  oa�pi�N   b�1   �E  'F  ch  mB  h__f ��?  |^F  ��	  |�a  �E1   i�E  i p��   �BF  NG  j�E  � jF  �jF  �jF  �nB  ��   ��F  lB  I� p��n   kPD  ����  �(G  lgD  �� l^D  �� t��  }tD  ׹ ~�D  �A  ��   ��F  l�A  � l�A  � l�A  /�  ��A  ��	   �l�A  Z� l�A  Z� l�A  Z� l�A  ��    o��p��   p���  o�p�N   ��1   �
   �fG  ~G  �h  mB  m� q*��   ��1  0�
   ��G  �G  �h  mB  �� q:��   �D  "O�G   �4  ��  "P�G  �1  "Q�G  ��  "W�G   �4  �^  "X�G  �U  #=H   	5  ��   #>H  �B  #?H  ��  #E2H   5  �B   #F2H  �C  #G2H  �e  #H2H  �8  #I2H  ��  #J2H  �

  #X�H   5  ��  #Y�H  ��
  #Z�H  ��   #`�H  *5  ��  #f�H   55  ��  #g�H  ��  #h�H  ��  #n�H   @5  ��	  #o�H  ��  #p�H  �H  #vI   K5  �`  #wI  �w  #xI  �   #yI  �~  #TI   V5  �   #�TI  ��  #�TI  �  #�TI  ��   #�TI  ��  #�TI  ��	  #�TI  ��  #��I   a5  �  #��I  �  #��I  ��  #��I  ��  #��I   l5  ��  #��I  ��  #��I  ��  #��I  �m  #�&J   w5  �	  #�&J  �2	  #�&J  ��  #�&J  �9  #�&J  �[  #�lJ   �5  �J  #�lJ  ��  #�lJ  �7  #�lJ  ��  #��J   �5  �I	  #��J  �$	  #��J  ��   #��J   �5  �N  #��J  �p  #��J   �5  ��  #��J  �:  #��J  ��  #��J  �d   #��J  ��  #�6K   �5  �  #�6K  ��  #�6K  ��	  #�bK   �5  ��  #�bK  �  #؁K   �5  ��  #فK  ��  #ځK  ��  #ہK  �+  #�K   �5  ��  #�K  ��   #�K  �  #��K   �5  ��
  #��K  ��  #��K  �  #�L   �5  �   #�L  �F  #�L  ��  #�>L   �5  ��  #�>L  ��  #�>L  ��  $3jL   6  ��  $4jL  ��   $8�L   6  ��  $9�L  �l	  $=�L  6  �N  $>�L  �^  $?�L  �L  $@�L  �a  $D�L  )6  �B  $E�L  ��	  $F�L  �  $G�L  �  $H�L  �y  $I�L  ��  % 4M   46  ��  %!4M  �1  .��  ��  ��  ��  ��  �   �  �  �!  �,  �8  �D  �P  �\  �h  �t  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  ��  �  �  ��  �Q  ���  �	Q�  �>  Y  .N  �4   ��  �1  �4    5   �M  � � �V  ح      ��  (  �  �  �  E   �  �  o  �	  �  qW  !s   int   "�   �  #  .  <h   `  Ds   �  Wh   �  _z   �  es   t   ms   a  us     ~s   �  �s   3  �s   �  �s   H  �s   y  �s     �s   s  �s   T   �s   �  �s   F  �s   �  �s   �  �s     �s   V  �s   3   �  s  N:   �  V:   \	  2s   o  7s   �  <s   �  Cs   �  s   �  3   	pO qO 	!�  std    	
@�  	5  	6.  	7H  
%  0�=  ��  �b  �3   Fe  �s   �3  �=  g  �  �   7  eq �<-  �  �  �  �   lt ��1  �  �  �  �   ��  eF  s   �  �  �  �   �K  �9  �  �  �   �(  
!  �    �  �  �   1  �A  �  ,  �  �  �   �5  �'  �  P  �  �  �   �3  �A  �  t  �  �  7   +  :  7  �  �   B  �C   �P  B  �  �   �B  $6  �  �  �  �   eof (�:  B  ?  ,N0  B  �    _� �,   �?  �%   �M  �  �* �e  �  +  1  �   �b  �3   �* �_e  �  V  \  �   \b  (a  q  |    �   �-  �  �  �  �  �   �-  P  �  �  �  �   � !4  �  �    s    cb  �Pc  �  �    s    �a  R(b           Fe  �B  �S  �YH    >  I    1   �c  <�c    b  h     �W  �B  �  �  �    �	  �   1  !a  *�a    �  �     !T  3   �E  +   	  �>  b�  �U  %7  �  �      �	   �   �  8.  �{  �   ]�  �  \�   �  �D  !�  �3  "�  U>  #�  &�  $�  �  %�  �*  &�   ڡ  '3   $�U  (3   %TL  )3   &�I  *3   'Q  +3   (�C  ,3   )�J  -3   *1  .�  ,o(  /3   0�U  03   1PL  13   2�I  23   3Q  33   4�C  43   5�J  53   6 )%  K�  H  s   �   GT  PS    $   'z  
�  $	,�  	-�   �� �� �� 2*  7�  8$   7  g  �  g  7  �    1  �     �  �  !h  �   �   =      !h  �   	   \  #  9  !h  9  "__n �      |  L  V  !h  �    �  d  n  !h  �    �  |  �  !h  9  "__n !s     �  �  �  !h  9  "__n �s    #t  �  "__c �   �  #�  �  "__c  �   �   �  �  	  !h  9  $%�&  T     %  "	  F	  !h  9  "__c �1  $%�&  �     I  T	  l	  !h  9  $%�&  >    #�  �	  &hR  $�	  &mR  $�	   �  �  '�  �   h  �	  �	  !h  9  "__s ��	  "__n ��    �  �	  �	  !h  9  $%�&  ,    �  (�  @�  ��  )�3  %  � )�D  &  �)Z*  &�  �* �  +�&  )�  �� ,__c +B  � -�  Y�0�  +�
  .�  +� /Y�   �
  0	  1�  b�   V.�  l�   *8�  2�  S*8�  3	  P   *P�  ,__n .�  � /}�   G  +� 1�  �� 4�	  }�   1$  .�	  �� .�	  λ .�	  �  5  ��   2.#  �� .,  ��   -�	  ��p�  DZ  .�	  � *p�  6�	  %� 7�  ����  /�  .�  G� /��   �  .�  Z� 8��   6	  m�   8��   0	  1�  ��   V.�  ��    9F	  ����  ..T	  � /��
   1  6^	  �� 1�  ��   B:�  .�  ��   8 �	   .T	  �� 8 �	   6^	  ��      ;	  ����  =.+	  ͼ ."	  � /��   �  68	  	� 1n  ��
   �:|  .�  �   8��   .+	  0� ."	  C� 8��   68	  	� 1�  ��   �.�  V�        �	  <U  =   �   <�   >  <B  ?  <�  E8   �   <B   F8  <C  G8  <e  H8  <8  I8  <�  J8  <

  X�   �   <�  Y�  <�
  Z�  =�   `�  �   <�  f�   �   <�  g�  <�  h�  <�  n�   �   <�	  o�  <�  p�  <H  v   �   <`  w  <w  x  <   y  <~  F   �   <   �F  <�  �F  <  �F  <�   �F  <�  �F  <�	  �F  <�  ��   �   <  ��  <  ��  <�  ��  <�  ��   �   <�  ��  <�  ��  <�  ��  <m  �	     <	  �	  <2	  �	  <�  �	  <9  �	  <[  �J     <J  �J  <�  �J  <7  �J  <�  �     <I	  �  <$	  �  <�   ��   "  <N  ��  <p  ��   -  <�  ��  <:  ��  <�  ��  <d   ��  <�  �   8  <  �  <�  �  <�	  �/   C  <�  �/  <  �L   N  <�  �L  <�  �L  <�  �L  <+  �   Y  <�  �  <�   �  <  �   d  <�
  �  <�  �  <  ��   o  <   ��  <F  ��  <�  ��   z  <�  ��  <�  ��  <D  O%   �  <�  P%  <1  Q%  <�  WN   �  <^  XN  <�  3k   �  <�  4k  <�   8�   �  <�  9�  <l	  =�  �  <N  >�  <^  ?�  <L  @�  <a  D�  �  <B  E�  <�	  F�  <  G�  <  H�  <y  I�  <�   '   �  <�  !'   Ǜ   Q  � �$ �V  ��      0�  �  (  �  �  �  L   �  �  o  �	  �  qW  !z   int   "%   #  .  <o   `  Dz   �  Wo   �  _�   �  ez   t   mz   a  uz     ~z   �  �z   3  �z   �  �z   H  �z   y  �z     �z   s  �z   T   �z   �  �z   F  �z   �  �z   �  �z     �z   V  �z   :   �  s  NA   �  VA   \	  2z   o  7z   �  <z   �  Cz   �  z   �  �  :   	pO qO !�  
std % W,  @�  ++ S��  Y�$ _;       ��  cN  (    �  ga  ;    %  0�=  �F  �b  �:   Fe  �z   �#  �F  �&  �  �3  �=  �  �2  �2   t  eq �<-  �2  �  �2  �2   lt ��1  �2  �  �2  �2   ��  eF  z     �2  �2  �   �K  �9  �  7  �2   �(  
!  �2  [  �2  �  �2   1  �A  �2    �2  �2  �   �5  �'  �2  �  �2  �2  �   �3  �A  �2  �  �2  �  t   +  :  t  �  �2     �C   �P       �2   �B  $6  �2    �2  �2   eof (�:    ?  ,N0    �2    E  
�Q  9Q  
p�  G0  
s�   �T  
t�  %  
{�  �  @5   %  
��  �  @5  �   �:  
�b;  �  �  �  F5   �T  
�4>  �  �  @5  �   �T  
�QM  �  �    F5   �F  
��?  L5    $  @5  �    I  
�O  L5  <  G  @5  �   (*  
�	H  Q  _  j  F5  �   �O  
�eT  Q  �  �  F5  �   �O  
́?  �  �  �  F5  R5   �$  �   �:  
Z�   _� �3   5�2  64  784  �?  �,   K  \p  w,   �e  _�  �4  cT4  �J  dZ4  ��  q7  =  r4   ��  sM  X  r4  x4   W  yd  r4  z     �  �J  p�   �B  �  �   !%  �   "�B  �  �  �4  �  x4   #�B  �  �4  z     �e  y  $[V  �  �  !�G  !�   <  x�  �4  {  �J  |  �J  .  `S  �,0  ~J  ��  �J  ��  �%  ��  �K  ��   I  ��  :!  �I4   %H  �:	  U   %�3  2�  %�G  7�  %t3  B�4  &�'  ��O  �4  'V  ��N  �2  �  �  �4   '3  �o+  �2  �    �4   (�P  ��O      �4   (�M  ��P  .  4  �4   (�,  �-  G  R  �4  �   '�+  ��R  �  i  o  �4   '3  �   �  �  �  �4  x4  x4   �/  !�B  �4  �  �  �  x4   (�O  �|6  �  �  �4  x4   )(  ��6  �  �  �4  x4   *�   �-  �  	  	  �4   +�1  o�*  �  )	  �4  x4  �    *�A  $n%  �  R	  X	  �4   *�A  (�I  �  p	  {	  �4  �   *"A  ,�%  �4  �	  �	  �4   *�1  2E)  %  �	  �	  �4   *�/  6;&  %  �	  �	  �4   )�>  :�>  �	  �	  �4   *S  A:2  �  
  
  �4  �  �   )�#  K�(  +
  @
  �4  �  �  �   *9  S>$  �  X
  h
  �4  �  �   *-U  [�7  �2  �
  �
  �4  �   ,�5  d�-  �
  �  �  �   ,	1  m�P  �
  �  �  �   ,�3  v\-  �
  �  �  :    ,nU  ��-    �  %  %   ,nU  �nG  +  �  1  1   ,nU  ��   K  �  �  �   ,nU  �IP  k  �  �  �   �J  �rR  z   �  �  �   )�=  ��H  �  �  �4  �  �  �   )V  �)  �  �  �4   -�'  �D*  �4  .�0  ��  �  �4   /�0  �    �4  x4   �0  �  *  �4  �4   �0  �:  O  �4  �4  �  �   �0  �_  y  �4  �4  �  �  x4   �0  ��  �  �4  �  �  x4   �0  ��  �  �4  �  x4   �0  ��  �  �4  �  :   x4   .�0  "�  �  �4  z    0�  *,Q  �4    #  �4  �4   0�  2�G  �4  <  G  �4  �   0�  =�%  �4  `  k  �4  :    0S� f�&  %  �  �  �4   0S� q�>  1  �  �  �4   1end y<  %  �  �  �4   1end �6;  1  �  �  �4   0I ��$  I       �4   0I ��7  =    %  �4   0��  �lC  I  >  D  �4   0��  �CM  =  ]  c  �4   0r ��R  �  |  �  �4   0�K  �r5  �  �  �  �4   0�3  �j=  �  �  �  �4   2�� �  �  �  �4  �  :    2�� ��F  �    �4  �   0I  v  �    $  �4   2�E  �|U  9  D  �4  �   2�1  -�  Y  _  �4   0�� 5�?  �2  x  ~  �4   0�:  D�6    �  �  �4  �   0�:  UW    �  �  �4  �   1at k
/    �  �  �4  �   1at ��7        �4  �   0�F  ��/  �4  %  0  �4  �4   0�F  �k:  �4  I  T  �4  �   0�F  ��H  �4  m  x  �4  :    0@  DA:  �4  �  �  �4  �4   0@  U�1  �4  �  �  �4  �4  �  �   0@  )�D  �4  �  �  �4  �  �   0@  ��*  �4      �4  �   0@  �6  �4  0  @  �4  �  :    2�G  -aN  U  `  �4  :    �3  �b*  �4  x  �  �4  �4   0�3  ^ 2  �4  �  �  �4  �4  �  �   0�3  �=  �4  �  �  �4  �  �   0�3  z�T  �4  �  �  �4  �   0�3  � @  �4    '  �4  �  :    2� ��E  <  Q  �4  %  �  :    0� �\+  �4  j  z  �4  �  �4   0� �u>  �4  �  �  �4  �  �4  �  �   0� g|=  �4  �  �  �4  �  �  �   0� "�@  �4  �    �4  �  �   0� 9k<  �4    2  �4  �  �  :    0� K�'  %  K  [  �4  %  :    0bL  d�R  �4  t  �  �4  �  �   0bL  t�2  %  �  �  �4  %   0bL  �L&  %  �  �  �4  %  %   0�%  �9F  �4  �  �  �4  �  �  �4   0�%  �|<  �4    7  �4  �  �  �4  �  �   0�%  ��T  �4  P  j  �4  �  �  �  �   0�%  ��A  �4  �  �  �4  �  �  �   0�%  b>  �4  �  �  �4  �  �  �  :    0�%  3%  �4  �  �  �4  %  %  �4   0�%  'V7  �4    ,  �4  %  %  �  �   0�%  <�+  �4  E  Z  �4  %  %  �   0�%  Q'S  �4  s  �  �4  %  %  �  :    0�%  vj.  �4  �  �  �4  %  %  �  �   0�%  ��9  �4  �  �  �4  %  %  �  �   0�%  �C  �4    &  �4  %  %  %  %   0�%  �>/  �4  ?  Y  �4  %  %  1  1   *�?  ��&  �4  q  �  �4  �  �  �  :    *�1  �O  �4  �  �  �4  �  �  �  �   ,)  �z-  �  �  �  :   x4   3+E  �3J  �    �  :   x4   0�5  ��)  �    2  �4  �  �  �   2n	 @D  G  R  �4  �4   0W�  �6  �  k  q  �4   0�A  %�A  �  �  �  �4   0��  ,Z5    �  �  �4   0�(  �;  �  �  �  �4  �  �  �   0�(  I�%  �  �    �4  �4  �   0�(  X�5  �    /  �4  �  �   0�(  �^   �  H  X  �4  :   �   0�(  v�S  �  q  �  �4  �4  �   0�(  	K  �  �  �  �4  �  �  �   0�(  �o?  �  �  �  �4  �  �   0�(  J5  �  �    �4  :   �   0NW  ��Q  �    *  �4  �4  �   0NW  /�I  �  C  X  �4  �  �  �   0NW  ��,  �  q  �  �4  �  �   0NW  ��;  �  �  �  �4  :   �   0�S  ��I  �  �  �  �4  �4  �   0�S  >T?  �  �    �4  �  �  �   0�S  05  �    *  �4  �  �   0�S  $S:  �  C  S  �4  :   �   0�>  2hL  �  l  |  �4  �4  �   0�>  SUB  �  �  �  �4  �  �  �   0�>  Q�2  �  �  �  �4  �  �   0�>  _�K  �  �  �  �4  :   �   0�4  qT  �    %  �4  �4  �   0�4  j�K  �  >  S  �4  �  �  �   0�4  ��5  �  l  |  �4  �  �   0�4  N.  �  �  �  �4  :   �   0U+  �)  u  �  �  �4  �  �   0��  �!1  z   �  �  �4  �4   0��  ��T  z        �4  �  �  �4   0��  ��O  z   9  X  �4  �  �  �4  �  �   0��  �;.  z   q  |  �4  �   0��  ��B  z   �  �  �4  �  �  �   0��  ��,  z   �  �  �4  �  �  �  �   �  3�) {$ �    ß  �  �  �  x4  (   E) ��* �  E  �  �  �  �  x4     �) ��$ �  r  �  �  �  �  x4   {* ��  �  f�  �  �4  �  �  x4   !T  :   4�E  h  4�F  �   5�&  5�7  u  6W  3Z  7�4  7�$  7q-  7c=  7o'  7�5   7�%  � 7�8  �7X)  �7�%  �7�  �7aO  �7Y=  � 7P  �� 7�C  ��7wS  �7�O  � 7�?  �7�5  �� 6
$ g�  7)W  7�   7�U  7�A  7�8  7�P   7EH  �� 6�4  ��  7O   7�7  7(  7�Q  7G  �� 6��  ��  7�R   7�-  7�1  7lO  �� 8b4 �   9�9  iZ  9�N  ��  �P  ��  :�4  $  
  ;dec $  :t-  $  ;hex $  :r'  $  :< $   ;oct $  @:� $  �<[)  $   <�%  "$   <�  &$   <dO  )$   <\=  ,$   <�P  /$    <�C  3$   @:zS  6$  �:�O  9$  J<�?  <$  9�  J�  :�7  N:      :(  Q:   :�Q  V:   :O  Y:    ;app lw   �  ;ate ow   ;in ww   ;out zw   ;cur ��   �  ;end ��    8�8  )!  .�  ��   �   8  z   �4   =�@  ]�   !  !  8  z   �4   !T  :   4�E  h   8�Y  �!  =�% g)!  G!  W!  <8  z   �4   .̾ ^h!  x!  <8  z   �4   !T  :   4�E  h   8�M  3#  0�-  P  �5  �!  �!  �5   �b  �:   0�* �e  �5  �!  �!  �5   0� � �5  �!  �!  �5   0�* �_e  �5  "  "  �5   0% ��" �5  5"  ;"  �5   2cb  �Pc  P"  ["  J6  z    0�-  �  �5  t"  z"  �5   2� !4  �"  �"  J6  z    =Z  ��!  �"  �"  J6  z    2��  �R�  �"  �"  J6  �5  �5  �5   2��  +�  �"  	#  J6  �5  �5   .�B �#   #  J6   !T  :   4�E  h   >8+ (@�!  A&  �!   ?�% S�   5# Nu  ?� VW#  $�b  D:   Fe  I  �#  J�  �&  K�  {'  M�!  �e  O�  /� b�#  �#  �4  �   /� o�#  �#  �4  �4  �   W#  @str ~n! W#  $  $  �4   Astr �� *$  5$  �4  �4   � �� I$  T$  �4  �   B��  ��& F&  3#  t$  z$  �4   B�[  �@ |#  	3#  �$  �$  �4   BZ  -�! |#  3#  �$  �$  �4  |#   BP� O( |#  3#  �$  �$  �4  |#   BY@ ��! �4  3#  %  &%  �4  �4  F&   B09  �� �#  3#  F%  [%  �4  �#  �  �   B=H  �} �#  3#  {%  �%  �4  �#  �   � �" �%  �%  �4  �4  �#  �#   �* �  �%  �%  �4   2� -! �%  �%  �4  �4  �4  �#   C� 3#  &  &  �4  z    �#  p#  �#  !T  :   4�E  h  4�F  �   3#  �>  
b�  D8 �)!  �'  )!   9�& 3#  !+ #i&  95# u  E�* 4�&  �&  �4  z   �4  �   E�* F�&  �&  �4  z   �4  �4  �   �&  F�* QQ&  �&  '  �4  z   �4   03F  \�* 5  %'  +'  
5   1str d& �&  D'  J'  
5   Gstr n _'  j'  �4  �4   !T  :   4�E  h  4�F  �   Q&  Dc  ���   �(  �    9�& �3#  !+ ��'  95# �u  E�% ��'  �'  5  z   �4  �   E�% �(  (  5  z   �4  5  �   �'  F�% ��'  6(  F(  5  z   �4   03F  �;' 5  _(  e(  "5   1str �� �'  ~(  �(  "5   Gstr ��& �(  �(  5  5   !T  :   4�E  h  4�F  �   �'  DS% ��)!  �)  �)   9�& 3#  !+ 	�(  95# u  E(% )  *)  (5  z   �4  �   E(% );)  U)  (5  z   �4  .5  �   �(  F'% 4�(  p)  �)  (5  z   �4   03F  ?� 45  �)  �)  :5   1str G� �(  �)  �)  :5   Gstr Q� �)  �)  (5  .5   !T  :   4�E  h  4�F  �   8$ ]*  Fk* ;�)  *  )*  ?L  z   �4   .l* >:*  J*  ?L  z   �4   !T  :   4�E  h   �(  Q  ד  ��*  �q  �N  ��  ��  � ��  �4  �T4  {�  �   �k  ��*  ��  ��  � ��  �4  �Z4  {�  �   �!  8�E  T+  F`V  �*  +  +  �7  z    .aV  � +  &+  �7   !T  :   4�E  h  Hi3 ~P4  H+  �7  J6    I*  sZ  n+  Z  Z   I�*  wZ  �+  Z  Z   I�% 	�S=  �+  J_Tp 3   S=  S=   Iͳ  	�S=  �+  J_Tp 3   S=  S=   I}�  ��2  �+  J_Tp :   x4  x4   IP* �s*  ,  8�  �  v5   I�% Z~*  7,  ��  �  �  �  N   K�% r~*  f�  �  �  �    L$   !��2  �  $,�  -�  K  :.  �e  =�  � ?�  "  @�  �4  AT4  �J  BZ4  �A  O�,  �,  `4   �A  Q�,  �,  `4  f4   �A  V -  -  `4  z    �
 Y51  �,  #-  .-  l4  �,   �
 ]�R  �,  F-  Q-  l4  �,   � c?  �,  i-  y-  `4  �,  �   _ m.   �-  �-  `4  �,  �,   �3  q89  �,  �-  �-  l4   .E  ��3  �-  �-  `4  �,  Z4   �(  ��(  �-  �-  `4  �,   J_Tp :    w,  MZD  �,0  NF�  ��   9��  �~*  9�4  ��*  9� ��*  .��  �`.  f.  p5   E��  �w.  �.  p5  v5   0*  ��}  5.  �.  �.  �5   0Ư  �?s  B.  �.  �.  �5   0�F  �Ϭ  �5  �.  �.  p5   0�F  ��  .  �.  /  p5  z    0a�  �
�  �5  /  "/  p5   0a�   ��  .  ;/  F/  p5  z    0�:  ,�  5.  _/  j/  �5  (.   0�F  		n  �5  �/  �/  p5  (.   0(*  ��  .  �/  �/  �5  (.   0 I  h�  �5  �/  �/  p5  (.   0�O  7k  .  �/  �/  �5  (.   0WC  ]�  v5  0  0  �5   {�  �  �  u   M8E  �K2  NF�  ��   9��  ��*  9�4  ��*  9� ��*  .��  �0  �0  X5   E��  ��0  �0  X5  ^5   0*  ���  T0  �0  �0  d5   0Ư  �p�  a0  �0  �0  d5   0�F  �5�  j5  �0  �0  X5   0�F  �÷  ,0  1  "1  X5  z    0a�  ��j  j5  ;1  A1  X5   0a�   �i  ,0  Z1  e1  X5  z    0�:  m�  T0  ~1  �1  d5  G0   0�F  	�u  j5  �1  �1  X5  G0   0(*  �  ,0  �1  �1  d5  G0   0 I  *�  j5  �1  �1  X5  G0   0�O  �  ,0  2  2  d5  G0   0WC  �i  ^5  22  82  d5   {�  �  �  u   ,0  .  OU  AI4  o2  �5  z    O9+  NI4  �2  �5  z    K;%  ��2  �  :   �    �� �� �� L2*  7�2  P8a   Qt  Q�  �  �  t  Q�  �  8"4  �{  "�   ]�  "�  \�  " �  �D  "!�  �3  ""�  U>  "#�  &�  "$�  �  "%�  �*  "&�   ڡ  "':   $�U  "(:   %TL  "):   &�I  "*:   'Q  "+:   (�C  ",:   )�J  "-:   *1  ".�  ,o(  "/:   0�U  "0:   1PL  "1:   2�I  "2:   3Q  "3:   4�C  "4:   5�J  "5:   6 I)%  "K�  84  z   �   RGT  "PC4  �2  �  # z   Q:   Q�  w,  Q.  .  �  Qp    z   �2  �  �  u  �  Q�  Q�  Qu  S3   �4  T �  �  3   3#  Q�#  A&  �#  p#  Q&  �  Q�&  i&  �'  �'  Q(  �'  �(  �(  QU)  �(  ]*  Q  b*  QQ  Qb*  ,0  Q�4  K2  Q,0  .  Q|5  �  P2  Q.  I4  UU2  �5  VXF  A�5  V\;  Az   WX�T  CI4    �!  �*  Y�!  �5  �5  Zh  �5   �5  Y�!  �5  6  Zh  �5   Y�!  6  6  Zh  �5   Y�!  (6  26  Zh  �5   Y"  @6  J6  Zh  �5   �!  Y;"  ^6  t6  Zh  t6  [__n �z    J6  Y�  �6  �6  Zh  �6   �4  Y["  �6  �6  Zh  �5   Yz"  �6  �6  Zh  t6  [__n !z    Y:	  �6  �6  Zh  �6   Y{	  �6  7  Zh  �6   Y�  7  7  Zh  7   �4  U�  77  W\__p ��    Y  E7  O7  Zh  O7   �4  Y�"  b7  u7  Zh  t6  Z#  �4   Uo2  �7  VXF  N�5  V\;  Nz    Y�  �7  �7  Zh  O7  ]__a �7   x4  Yc  �7  �7  Zh  �6   �*  Y�*  �7  �7  Zh  �7  Z#  �4   �7  �   Y�   8  28  Zh  28  Z#  �4  Z�!  78   8  �4  )!  Y2!  P8  l8  Zh  l8  Z#  �4  Z�!  q8   <8  �4  Y�   �8  �8  Zh  28  Z#  �4  Z�!  �8   �4  U�  �8  VhR  ��8  VmR  ��8   �2  �2  YR  �8  �8  Zh  O7   Y4  �8  9  Zh  O7  ]__n ��   Y  9  #9  Zh  �6   U�  D9  VhR  �D9  VmR  �I9   �2  �2  U  }9  ^�e  �2  ^�e  �2  [__n �   U�
  �9  [__d d�  [__s d�  [__n d�   U�  �9  [__c �9   �2  U�  �9  [__c  �9   �2  U   :  ^hR  $:  ^mR  $:   �2  �2  _  U/  .:  [__c ,.:   �2  UT+  T:  ]__a sZ  ]__b sZ   Y�"  b:  �:  Zh  t6  ^�  ��5  ^;�  ��5  ^P�  ��5   Y�%  �:  �:  Zh  �:  WX�
 �4    �4  Y�"  �:  �:  Zh  t6  ^M�  +�5  ^u�  +�5   Yq  �:  ;  Zh  �6   Un+  #;  ]__a wZ  ]__b wZ   YD  1;  ;;  Zh  ;;   �4  Y�  N;  c;  Zh  c;  VQ  
��   @5  Y�  v;  �;  Zh  �;   F5  Y�,  �;  �;  Zh  �;   `4  Y'  �;  �;  Zh  �;   r4  Y�,  �;  �;  Zh  �;  Z#  �4   YX  �;  <  Zh  �;  Z#  �4   Y�,  <  <  Zh  �;  <   f4  Y=  1<  F<  Zh  �;  ]__a sF<   x4  Y�  Y<  c<  Zh  �6   `�  t<  �<  Zh  �<  Z#  �4   �4  Y	#  �<  �<  Zh  t6   Y�  �<  �<  Zh  ;;  Z#  �4   Y+  �<  �<  Zh  �7   Y�  �<  =  Zh  �<  ^v�  �  [__a =   x4  _�  Y�  &=  0=  Zh  ;;   Y�#  >=  S=  Zh  �:  V^F  b�   Q�4  U�+  �=  J_Tp 3   ]__a 	ك=  ]__b 	و=   S=  S=  U�+  �=  J_Tp 3   ]__a 	·=  ]__b 	¼=   S=  S=  U�+  �=  J_Tp :   �=  �=   x4  x4  U�+  >  8�  �  >   v5  U,  6>  ��  �  Vz  Z�  V�l  Z�  N   U�2  U>  �  :   VŐ   ��   U7,  >  f�  �  Vz  r�  V�l  r�   U+  �>  [__p ��  ^۶  ��  ^nh  ��   U�   ?  ß  �  V�|  |�  V�h  |�  ]__a | ?  (  WX�  ��  \__r ��4    x4  U  C?  �  �  ^�|  ��  ^�h  ��  [__a �C?    a x4  UE  �?  �  �  ^�|  ��  ^�h  ��  [__a ��?  a x4  Yr  �?  �?  f�  �  Zh  ;;  V�|  �  V�h  �  ]__a ��?   x4  Y�  �?  �?  Zh  ;;  ^�^  *�?   �4  bT$  `�6   �@  �@  ch  �:  n� dd�2   e�&  �F&  �� f�:  p�   �g�:  Ž dp�   h�:  ٽ fT:  x�   �g�:  �� gw:  	� gk:   � gb:  7�      bz$  ��F   ��@  ZA  ch  �:  K� d��B   e�&  �|#  v� e�
 ��4  �� i�:  ���  �?A  g�:  �� j�  h�:  ׾ fT:  ��   �g�:  � gw:  � gk:  -� gb:  A�    f�9  ��   �g�9  T�    b�$  ��W   �qA  |B  ch  �:  v� k__c .|#  �� j �  e�&  0|#  ׿ j �  X �  5�4  l�   :B  X�# 8�4  e8 ;�4  � m#9  �   :�A  n-9  g89  9�  m�9  �   9B  g�9  N�  oP6  �8�  >g^6  f� gg6  z�   iP6  0�P�  F`B  g^6  �� gg6  ��  f:  3�   Gg!:  ��     p�7  ��"   ��B   C  g�7  �� g�7  �� iu7  ��h�  ��B  q�7  g7  � o�5  ��h�  Vq�5  g�5  � jh�  h�5  6�    rʀ�   s�%  @C  #C  Zh  �:  Z#  �4   t C  @ P�`   �>C  SD  uC  � i�<  Y���  @4D  g�<  V� v�6  Y���  #�C  g�6  V� w�6  Y�   -g�6  V�   x�7  e���  #g�7  �� g�7  �� d��    g�7  �� g�7   � iu7  ��Ю  �(D  q�7  g7  � o�5  ��Ю  Vq�5  g�5  � jЮ  h�5  (�    r���     fT7  m�   @gb7  H� y�  t C  ) ��`   �nD  �E  uC  � i C  ���  @�E  gC  g� i�<  �� �  @�E  g�<  �� v�6  �� �  #�D  g�6  �� w�6  ��   -g�6  ��   x�7  ��8�  #g�7  �� g�7  �� d��    g�7  � g�7  ;� iu7  ��P�  �tE  q�7  g7  N� o�5  ��P�  Vq�5  g�5  N� jP�  h�5  c�    r��     fT7  ��   @gb7  �� y��  r����   Y (  �E  �E  Zh  �E  Z#  �4  Z�!  �E   5  �4  t�E  F$ ��   ��E  FG  u�E  � v C  �h�  �*G  gC  �� i�<  ���  @G  g�<  �� v�6  ���  #qF  g�6  �� w�6  �   -g�6  ��   x�7  3�ȯ  #g�7  � g�7  3� dp�    g�7  Q� g�7  ~� iu7  p��  ��F  q�7  g7  �� o�5  p��  Vq�5  g�5  �� j�  h�5  ��    r���     oT7  ;���  @gb7  �� yQ�  x�7  H��  �n�7  y_�  Y�&  TG  pG  Zh  pG  Z#  �4  Z�!  uG   �4  �4  tFG  u ���   ��G  �H  uTG  � v C  ��(�  R�H  gC  �� i�<  ��P�  @�H  g�<  � v�6  ��p�  #H  g�6  � w�6  ��   -g�6  �   x�7  ����  #g�7  O� g�7  |� d�    g�7  �� g�7  �� iu7  ���  ��H  q�7  g7  �� o�5  ���  Vq�5  g�5  �� j��  h�5  ��    r+��     oT7  ����  @gb7  � y��  x�7  ��а  Rn�7  y��  t�E  �  P��   ��H  wJ  u�E  � v�E  Y��  �mJ  g�E  4� v C  Y� �  �MJ  gC  ^� i�<  Y� �  @.J  g�<  �� v�6  Y�@�  #�I  g�6  �� w�6  Y�   -g�6  ��   x�7  s�X�  #g�7  �� g�7  �� d��    g�7  � g�7  :� iu7  ��p�  �"J  q�7  g7  M� o�5  ��p�  Vq�5  g�5  M� jp�  h�5  b�    r���     fT7  {�   @gb7  �� y��  w�7  ��   �g�7  �� y��  r����   tFG  V( ���   ��J  L  uTG  � vFG  ����  RL  gTG  �� v C  ����  R�K  gC  � i�<  ����  @�K  g�<  @� v�6  ���  #(K  g�6  @� w�6  ��   -g�6  @�   x�7  ���  #g�7  r� g�7  �� dP�    g�7  �� g�7  �� iu7  P��  ��K  q�7  g7  �� o�5  P��  Vq�5  g�5  �� j�  h�5  �    rk��     fT7  �   @gb7  2� y.�  w�7  .�   Rg�7  W� y@�  rH���   YZ)  L  5L  Zh  5L  Z#  �4  Z�!  :L   (5  �4  �)  Y*  SL  oL  Zh  oL  Z#  �4  Z�!  tL   ?L  �4  tL  �( ���   ��L  �M  uL  � v C  ��(�  5�M  gC  �� i�<  ��P�  @�M  g�<  �� v�6  ��p�  #M  g�6  �� w�6  ��   -g�6  ��   x�7  ����  #g�7  �� g�7  %� d��    g�7  C� g�7  p� iu7  ����  ��M  q�7  g7  �� o�5  ����  Vq�5  g�5  �� j��  h�5  ��    r �     oT7  ����  @gb7  �� y��  x�7  ��в  5n�7  y��  tL  C# @ �   ��M  vO  uL  � vL  I �  5lO  gL  �� v C  I  �  5LO  gC  � i�<  I  �  @-O  g�<  9� v�6  I @�  #�N  g�6  9� w�6  I    -g�6  9�   x�7  j X�  #g�7  k� g�7  �� d�     g�7  �� g�7  �� iu7  � p�  �!O  q�7  g7  �� o�5  � p�  Vq�5  g�5  �� jp�  h�5  �    r� �     fT7  r    @gb7  +� y�   w�7  �    5g�7  P� y�   r� ��   t0=  �#  Z   ��O  P  u>=  � uG=  �m�<  9   c�O  g�<  �� yA f=  K   cg&=  �� w�<  K   �n =  g�<  �� g�<  ��    Y�#  P  1P  Zh  1P  WX�&  �W#  Wn�<     �4  tP  n! `�   �QP  �T  uP  �z��  �T  {P  � m=  n	   ��P  g&=  �� w�<  n	   �n =  g�<   � g�<  ��   i�?  ���  �{Q  g�?  L� g�?  y� g�?  �� g�?  �� iH?  ���  �WQ  gs?  L� gg?  y� g[?  �� j��  x?  ���  �g0?  L� g$?  y� g?  �� j��  r��>      f�<  �   �n =  n�<  g�<  ��   i�?  �г  ��Q  g�?  �� g�?  �� r�`   i�<  ��  ��R  g�<  � v�6  ��  #�Q  g�6  � w�6  �   -g�6  �   x�7  �(�  #g�7  #� g�7  E� d�    g�7  c� g�7  �� iu7  �@�  ��R  g�7  �� g7  �� o�5  �@�  Vg�5  �� g�5  �� j@�  h�5  ��    r��     i�?  �X�  �iS  g�?  �� g�?  '� g�?  :� g�?  N� iH?  �p�  �ES  gs?  �� gg?  '� g[?  :� jp�  x?  �p�  �g0?  �� g$?  '� g?  :� jp�  r��>      f�<  �   �n =  n�<  g�<  ��   i�?  ���  ��S  g�?  �� g�?  �� r�`   i�?   ��  ��S  g�?  �� g�?  � r`   m�<     �5T  g�<  � |�6     #T  g�6  �  w�7  "   #g�7  .� g�7  [� }1|B  ~Rus   d1   g�<  n� |�6  1   #eT  g�6  n�  w�7  6   #g�7  �� g�7  �� }E|B  ~Rut    rN��   t�:    PB   ��T  U  g�:  �� dW;   h�:  �� fT:  h(   �g�:   � gw:   � gk:   � gb:  3�    b�%  �T   �'U  �U  ch  �:  G� M�  �4  �u�  �4  ��Q  �#  r� v�:  ���  �U  u�:  �u�:  �g�:  ��  |�6  �   �U  g�6  �� g�6  ��  w�6  �   
g�6  �� g�6  �   b�%   �   ��U  �W  �h  �:  � ���  ��4  �k__i �#  /� �__o �#  �jд  e�
 �4  [� e8 �4  �� e�% ��4  �� e{# ��4  � m�7     �V  g�7  V� w�6     �g�6  V� w�6     -g�6  V�    i3:  �  ��V  �H:  g=:  ��  m9     � W  g9  ��  m3:      �$W  �H:  g=:  �  mT:  A   �\W  g�:  2� gw:  P� gk:  �� gb:  ��  mT:  w   ��W  g�:  � gw:  � gk:  � gb:  �  rwU  r�U    Y5$  �W  �W  Zh  �:  V^F  ��  WXR'  ��#    t�W  � �@   ��W  vX  u�W  � u�W  �j �  h�W  (� i�7  ��  �bX  g�7  j� w�6  �   �g�6  j� w�6  �   -g�6  j�    r��U  r��U    b�$  �@   ��X  Y  �h  �:  � �__s ��4  ��__n �F&  �i#;  0�  ��X  g1;  �� |�7     .�X  g�7  ��  r�   r'�U   Y@  Y  9Y  Zh  ;;  [__c -:   W�R'  /�    b�$  0�  �PY  �]  �h  �:  � �__c P|#  �zH�  �]  e8 R�4  �� X �  V�4  e� Z&  <� e5 [&  �� e�" \�4  �� X� b&  i9  Rp�  Z�Y  g9  ��  z��  �]  e�* n&  � XR'  p&  �Y�  qW#  �\mY=  �   o4Z  nw=  nl=   m=  �   qyZ  g&=  ;� w�<  �   �n =  g�<  s� g�<  ;�   iY  ���  u�[  gY  �� gY  �� j��  h*Y  �� |�7  �   /�Z  g�7  �� w�6  �   �g�6  �� w�6  �   -g�6  ��    |�8     2%[  g�8  �� g�8  %�  |�6     3][  g�6  =� w�6     -g�6  =�   v�8  ��  3�[  g�8  _� g�8  � d�   g�8  �� g�8  �� m77  �   շ[  nE7   f�8  �   �n�8  g�8  ��    r�$    i�<  =ص  x�\  g�<  �� v�6  =�  #6\  g�6  �� w�6  =   -g�6  ��   w�7  F:   #g�7  �� g�7  %� dR.   g�7  8� g�7  e� iu7  R�  ��\  g�7  x� g7  �� o�5  R�  Vg�5  x� g�5  �� j�  h�5  ��    rp�     m�=  �    p�\  g�=  �� g�=  ��  m�<  �   xj]  u�<  ud�|�6  �   #6]  u�6  ud� w�7  �   #g�7  � g�7  ?� }�|B  ~Ruc   r�$  r��  r#2  r=�U   m�6  |   |�]  g�6  R� g�6  e�  f:  �   Xn!:    r���   Y$  �]  �]  Zh  �:  ]__s ��]   �4  t�]  �  ;   �^  _  u�]  � u�]  �i�7   �  �y^  g�7  y� x�6  8�  �g�6  y� x�6  P�  -g�6  y�    m�W     �_  g�W  �� g�W  �� d   h�W  �� i�7  $h�  �_  g�7  �� w�6  $   �g�6  �� w�6  $   -g�6  ��    r6�U    r�   Y�#  $_  D_  Zh  �:  V�^  oD_  V^F  p�   �4  t_  �) @�   �d_  a  u$_  � u-_  �u8_  �m�<  O9   q�_  g�<  �� y� i�7  ���  q�_  g�7  5� x�6  ���  �g�6  5� x�6  ���  -g�6  5�    i�W  �ȶ  r~`  g�W  l� g�W  �� jȶ  h�W  �� i�7  ��  �s`  g�7  � w�6  �   �g�6  � w�6  �   -g�6  �    r��U    m�<  �   q�`  g�<  0� |�6  �   #�`  g�6  0�  w�7  �   #g�7  E� g�7  r� }�|B  ~Rug   mT7  �   qa  ub7  Sy y�r��   b&%   E  �2a  �b  �h  �:  ��Q  ��#  ��@  ��  ��^F  ��  �j��  ��&  ��#  � e�
 ��2  �� e8 ��2  0� eK( ��4  e� e�|  ��b  �� i3:  7 �  ��a  gH:  �� �=:   i@;  =@�  �b  qW;  uN;  �  m3:  `   �'b  gH:  �� �=:   jX�  e�% ��#  � e� ��#  �� i�:  �p�  ��b  g�:  �� jp�  h�:  � oT:  ���  �g�:  t� gw:  t� gk:  t� gb:  ��    mT:  *   ��b  g�:  �� gw:  �� gk:  �� gb:  ��  rkU     &  b[%  p	  �c  �d  �h  �:  ��j(  ň#  � �^F  ��  �j��  ��&  ǈ#  � e�
 Ȋ4  D� e8 Ɋ4  X� e�|  ��b  l� i3:  �	��  ȝc  gH:  �� �=:   m@;  �	   ��c  qW;  gN;  ��  m3:  �	   ��c  gH:  �� �=:   jط  X%  � &  e� ъ4  !� i�:  �	�  �cd  g�:  A� j�  h�:  w� oT:  
�  �g�:  �� gw:  �� gk:  �� gb:  ��    mT:  j
   ֛d  g�:  �� gw:  �� gk:  � gb:  3�  r�
U     YW!  �d  �d  Zh  l8  Z#  �4  Z�!  �d   �4  Y�&  �d  e  Zh  pG  Z#  �4  Z�!  e  ^^F  4�   �4  t�d  ]) �
�   �,e  `f  u�d  � u�d  �u�d  �v�d  �
 �  5te  g�d  F� g�d  �� r�
8+   v0=  �
8�  5�e  gG=  �� g>=  �� i�<  �
X�  c�e  g�<  �� y f=     cg&=  4� w�<     �n =  g�<  v� g�<  4�    v;  p�  5#f  �;  g;  ��  |B8  K   5Hf  ub8  v�uP8  S r48+  yKrb��   t�d  � p  �{f  �g  u�d  � u�d  �|�<  |I   5�f  g�<  �� y� |�d  �   5�f  u�d  �	�g�d  � r�8+   v0=  ���  5kg  gG=  7� g>=  o� i�<  ���  c)g  g�<  o� y/ f=  9   cg&=  �� w�<  9   �n =  g�<  � g�<  ��    v;  /��  5�g  g;  *� g;  J�  |�7  p   5�g  u�7  s0�y� rO8+  yjr���   Y�&  �g  h  Zh  pG  Z#  �4  Z�!  h  ^�^  Fh  ^^F  G�   �4  �4  t�g  �" �K  �4h  �j  u�g  � u�g  �u�g  �uh  �v�d  �ظ  H�h  g�d  v� g�d  �� r�8+   v_  ��  HOj  g8_  �� g-_  a� g$_  �� i�<  � �  q�h  g�<  �� y i�7  H�  q&i  g�7  � x�6  `�  �g�6  � x�6  x�  -g�6  �    m�W  C    r�i  g�W  J� g�W  �� dC    h�W  �� i�7  O��  ��i  g�7  � w�6  O   �g�6  � w�6  O   -g�6  �    ra�U    m�<  �   q'j  g�<  ,� |�6  �   #�i  g�6  ,�  w�7  �   #g�7  A� g�7  n� }�|B  ~Rug   mT7  �   qIj  gb7  �� y� y@ v;  ���  Htj  �;  g;  ��  |B8  �   H�j  gb8  �� gP8  ��  rq8+  r���  y� t�g  �' ��  ��j  im  u�g  � u�g  �uh  �|�<  �I   H	k  g�<  �� y� |�d  5   H<k  u�d  �	�g�d  5� rS8+   v;  Sȹ  Hck  g;  k� g;  ��  v_  V�  H.m  g8_  �� g-_  X� g$_  �� i�<  V �  q�k  g�<  �� y� i�7  �P�  ql  g�7  #� x�6  �h�  �g�6  #� x�6  ���  -g�6  #�    m�W  �    r�l  g�W  [� g�W  �� d�    h�W  :� i�7  ���  ��l  g�7  Y� w�6  �   �g�6  Y� w�6  �   -g�6  Y�    r��U    m�<     qm  g�<  n� |�6     #�l  g�6  n�  w�7     #g�7  �� g�7  �� }%|B  ~Rug   mT7  %   q(m  gb7  �� y7 y� |�7  :   HQm  g�7  �� yJ r�8+  rR��  y[ tFG  v& p�   ��m  �n  uTG  � ufG  �v C  ���  R�n  gC  �� i�<  �Ⱥ  @�n  g�<  � v�6  ��  #n  g�6  � w�6  �   -g�6  �   x�7  � �  #g�7  Q� g�7  ~� d�    g�7  �� g�7  �� iu7  ��  ��n  q�7  g7  �� o�5  ��  Vq�5  g�5  �� j�  h�5  ��    r��     fT7  �   @gb7  � y�  wB8  �   Rgb8  6� gP8  [�   b'  �   ��n  o  �h  o  �  
5  b+'   �   �#o  �s  �h  o  �vP  0�  e�s  gP  z� j0�  �P  m=  	   ��o  g&=  �� w�<  	   �n =  g�<  � g�<  ��   i�?  &H�  �hp  g�?  1� g�?  ^� g�?  q� g�?  �� iH?  &`�  �Dp  gs?  1� gg?  ^� g[?  q� j`�  x?  &`�  �g0?  1� g$?  ^� g?  q� j`�  r5�>      f�<  6   �n =  n�<  g�<  ��   i�?  9x�  ��p  g�?  �� g�?  �� rD`   i�<  D��  ��q  g�<  �� v�6  D��  #�p  g�6  �� w�6  D   -g�6  ��   x�7  Mл  #g�7  � g�7  *� d�    g�7  H� g�7  u� iu7  ��  �q  g�7  �� g7  �� o�5  ��  Vg�5  �� g�5  �� j�  h�5  ��    r��     i�?  ` �  �Vr  g�?  �� g�?  � g�?  � g�?  3� iH?  `�  �2r  gs?  �� gg?  � g[?  � j�  x?  `�  �g0?  �� g$?  � g?  � j�  ro�>      f�<  p   �n =  n�<  g�<  m�   i�?  s0�  ��r  g�?  m� g�?  �� r~`   i�?  �H�  ��r  g�?  �� g�?  �� r�`   m�<  �   �"s  g�<  �� |�6  �   #�r  g�6  ��  w�7  �   #g�7  � g�7  @� }�|B  ~Rus   d�   g�<  S� |�6  �   #Rs  g�6  S�  w�7  �   #g�7  g� g�7  �� }�|B  ~Rut     r���   bJ'  �@   ��s  �t  �h  pG  � �__s n�t  �x�]  �`�  ou�]  �g�]  �� i�7  ���  �5t  u�7  �x�6  ���  �u�6  �x�6  ���  -u�6  �   m�W     ��t  g�W  �� g�W  �� d   h�W  � i�7  ȼ  ��t  g�7   � w�6     �g�6   � w�6     -g�6   �    r*�U    r�    �4  Y�'  �t  u  Zh  �E  Z#  �4  Z�!  u  ^^F  ��   �4  t�t  y' 0�   �.u  bv  u�t  � u�t  �uu  �v8  ?�  �vu  g(8  5� g8  w� rY8+   v0=  B��  � v  gG=  �� g>=  �� i�<  B�  c�u  g�<  �� y� f=  �   cg&=  #� w�<  �   �n =  g�<  e� g�<  #�    v;  �0�  �%v  �;  g;  y�  |v8  �   �Jv  u�8  v�u�8  S r�8+  y�r���   t�t  �(    �}v  �w  u�t  � uu  �|�<  I   ��v  g�<  �� y |8  U   ��v  n(8  g8  �� rl8+   v0=  lH�  �fw  gG=  &� g>=  ^� i�<  lh�  c$w  g�<  ^� y� f=  �   cg&=  �� w�<  �   �n =  g�<  � g�<  ��    v;  ���  ��w  g;  � g;  9�  |�7  �   ��w  u�7  s,�y	 r�8+  y�r��   Y�'  �w  
x  Zh  �E  Z#  �4  Z�!  
x  ^�^  �x  ^^F  ��   �4  5  t�w  *  @  �/x  �z  u�w  � u�w  �u�w  �u�w  �v8  /��  �x  g(8  e� g8  �� rI8+   v_  K��  �Jz  g8_  �� g-_  P� g$_  �� i�<  K�  q�x  g�<  �� y� i�7  ��  q!y  g�7  �� x�6  � �  �g�6  �� x�6  �8�  -g�6  ��    m�W  �    r�y  g�W  9� g�W  �� d�    h�W  �� i�7  �P�  ��y  g�7  � w�6  �   �g�6  � w�6  �   -g�6  �    r��U    m�<     q"z  g�<  � |�6     #�y  g�6  �  w�7     #g�7  0� g�7  ]� }!|B  ~Rug   mT7  !   qDz  gb7  p� y3 y� v;  \h�  �oz  �;  g;  ��  |v8  8   ��z  g�8  �� g�8  ��  r�8+  rO��  yX t�w  5 `�  ��z  ]}  u�w  � u�w  �u�w  �|�<  lI   �{  g�<  �� yu |8  �   �0{  n(8  g8  $� r�8+   v;  ���  �W{  g;  Z� g;  ��  v_  ���  �"}  g8_  �� g-_  G� g$_  � i�<  ��  q�{  g�<  � y$ i�7  $�  q�{  g�7  � x�6  $(�  �g�6  � x�6  $@�  -g�6  �    m�W  N    r�|  g�W  J� g�W  �� dN    h�W  )� i�7  ZX�  ��|  g�7  H� w�6  Z   �g�6  H� w�6  Z   -g�6  H�    rl�U    m�<  �   q�|  g�<  ]� |�6  �   #�|  g�6  ]�  w�7  �   #g�7  r� g�7  �� }�|B  ~Rug   mT7  �   q}  gb7  �� y� yK |�7  �   �E}  g�7  �� y� ru8+  r���  y� t�E  =& ��   �x}  �~  u�E  � u�E  �v C  p�  ��~  gC  �� i�<  ��  @�~  g�<  � v�6  ��  #�}  g�6  � w�6     -g�6  �   x�7  ��  #g�7  @� g�7  m� dP    g�7  �� g�7  �� iu7  Pؿ  ��~  q�7  g7  �� o�5  Pؿ  Vq�5  g�5  �� jؿ  h�5  ��    rk�     fT7      @gb7   � y3  wv8  3   �g�8  %� g�8  J�   bF(  p   ��~  �~  �h  �~  �  "5  be(  ��   �  ��  �h  �~  �vP  ��  �|�  gP  i� j�  �P  m=  �	   ��  g&=  �� w�<  �	   �n =  g�<  �� g�<  ��   i�?  ��  �\�  g�?     g�?  M  g�?  `  g�?  t  iH?  � �  �8�  gs?     gg?  M  g[?  `  j �  x?  � �  �g0?     g$?  M  g?  `  j �  r��>      f�<  �   �n =  n�<  g�<  �    i�?  �8�  ���  g�?  �  g�?  �  r�`   i�<  �X�  ��  g�<  �  v�6  �x�  #߀  g�6  �  w�6  �   -g�6  �    x�7  ���  #g�7  �  g�7   d     g�7  7 g�7  d iu7   ��  �s�  g�7  w g7  � o�5   ��  Vg�5  w g�5  � j��  h�5  �    r�     i�?  ���  �J�  g�?  � g�?  � g�?   g�?  " iH?  ���  �&�  gs?  � gg?  � g[?   j��  x?  ���  �g0?  � g$?  � g?   j��  r��>      f�<  �   �n =  n�<  g�<  \   i�?  ���  �y�  g�?  \ g�?  � r�`   i�?   �  ���  g�?  � g�?  � r-`   m�<  <   ��  g�<  � |�6  <   #�  g�6  �  w�7  B   #g�7   g�7  / }Q|B  ~Rus   dQ   g�<  B |�6  Q   #F�  g�6  B  w�7  V   #g�7  V g�7  � }e|B  ~Rut     rn��   b�(  p@   ���  Ǆ  �h  �E  � �__s �Ǆ  �x�]  u �  �u�]  �g�]  � i�7  u@�  �)�  u�7  �x�6  uX�  �u�6  �x�6  up�  -u�6  �   m�W  �   ���  g�W  � g�W  � d�   h�W  � i�7  ���  ���  g�7   w�6  �   �g�6   w�6  �   -g�6      r��U    r��    5  Y)*  ڄ  ��  Zh  oL  Z#  �4  Z�!  ��   �4  Y)  	�  1�  Zh  5L  Z#  �4  Z�!  1�  [__m �   �4  t��  �  �  �Q�  Æ  u	�  � u�  �u$�  �v̄  ���  �  g�  $ gڄ  v |�d  �"   ?��  g�d  � g�d  v r�8+   |8  �   ?�  g(8  � g8  P r�8+   wB8  �   ?gb8  � gP8  �   v0=   ��  ��  gG=  � g>=  � i�<   ��  c[�  g�<  � yc f=  m   cg&=  ; w�<  m   �n =  g�<  � g�<  ;    r�8+  r���  y�y�r���   t��  �# �A  �ކ  Z�  u	�  � u$�  �|�<  �I   �  g�<  � y� |̄  %6   ��  g�  � gڄ  ) |�d  %    ?c�  n�d  g�d  ) rC8+   w8  E   ?g(8  _ g8  � r[8+    v0=  [ �  �  gG=  � g>=  � i�<  [�  c؇  g�<  � y� f=  �   cg&=  M w�<  �   �n =  g�<  � g�<  M    |�7  �   =�  u�7  s4�y	 r�8+  y�y�r��   Y*)  h�  ��  Zh  5L  Z#  �4  Z�!  ��  ^�^  )��  [__m *�   �4  .5  tZ�  ]"  �  ���  x�  uh�  � uz�  �u��  �u��  �v̄  /0�  +��  g�  � gڄ  
	 |�d  /"   ?7�  g�d  @	 g�d  
	 rQ8+   |8  Q   ?g�  g(8  �	 g8  �	 rm8+   wB8  �    ?gb8  :
 gP8  O
   v_  �P�  +R�  g8_  b
 g-_  �
 g$_  �
 i�<  �p�  q܉  g�<  �
 y� i�7  ���  q-�  g�7  r x�6  ���  �g�6  r x�6  ���  -g�6  r    i�W  ���  r��  g�W  � g�W   j��  h�W  � m�7  
   ���  g�7  � w�6  
   �g�6  � w�6  
   -g�6  �    r�U    m�<  M   q*�  g�<  � |�6  M   #��  g�6  �  w�7  S   #g�7  � g�7   }b|B  ~Rug   mT7  b   qL�  gb7    yt y� r*8+  y�r���  r���  y� tZ�  I ��  ���  T�  uh�  � u��  �u��  �|�<  �I   +΋  g�<  5 y� |̄  6   +M�  g�  � gڄ  � |�d      ? �  n�d  g�d  � r38+   w8  5   ?g(8  � g8  . rK8+    v_  K��  +�  g8_  � g-_  � g$_   i�<  K�  q��  g�<   y� i�7  �8�  q�  g�7  � x�6  �P�  �g�6  � x�6  �h�  -g�6  �    i�W  ���  r~�  g�W  � g�W  - j��  h�W  � i�7  ���  �s�  g�7  � w�6  �   �g�6  � w�6  �   -g�6  �    r��U    m�<     q�  g�<  � |�6     #��  g�6  �  w�7     #g�7  � g�7  * }!|B  ~Rug   mT7  !   q�  gb7  = y3 y� |�7  F!   +7�  g�7  R yV r�8+  yCr^��  yp tL  }+ ��   �o�  �  uL  � u+L  �v C  ���  5��  gC  g i�<  ���  @��  g�<  � |�6  �   #��  g�6  � w�6  �   -g�6  �   x�7  ���  #g�7  � g�7  � d    g�7   g�7  C iu7  �  �~�  q�7  g7  V o�5  �  Vq�5  g�5  V j�  h�5  k    r+�     fT7  �   @gb7  � y�  wEL  �2   5geL  � gSL  � |v8  �   ;�  g�8  � g�8    wB8  �   ;gb8  > gP8  c    b�)  0   �.�  <�  �h  <�  �  :5  b�)  @�   �X�  ǔ  �h  <�  �vP  N �  H��  gP  � j �  �P  m=  N	   �Ґ  g&=  � w�<  N	   �n =  g�<   g�<  �   i�?  f8�  ���  g�?  9 g�?  f g�?  y g�?  � iH?  fP�  �y�  gs?  9 gg?  f g[?  y jP�  x?  fP�  �g0?  9 g$?  f g?  y jP�  ru�>      f�<  v   �n =  n�<  g�<  �   i�?  yh�  �̑  g�?  � g�?  � r�`   i�<  ���  ���  g�<  � v�6  ���  # �  g�6  � w�6  �   -g�6  �   x�7  ���  #g�7   g�7  2 d�    g�7  P g�7  } iu7  ���  ���  g�7  � g7  � o�5  ���  Vg�5  � g�5  � j��  h�5  �    r��     i�?  ���  ���  g�?  � g�?   g�?  ' g�?  ; iH?  ��  �g�  gs?  � gg?   g[?  ' j�  x?  ��  �g0?  � g$?   g?  ' j�  r��>      f�<  �   �n =  n�<  g�<  u   i�?  � �  ���  g�?  u g�?  � r�`   i�?  �8�  ��  g�?  � g�?  � r�`   m�<  �   �W�  g�<   |�6  �   ##�  g�6    w�7     #g�7   g�7  H }|B  ~Rus   d   g�<  [ |�6     #��  g�6  [  w�7     #g�7  o g�7  � }%|B  ~Rut     r.��   b�)  0@   �ޔ  �  �h  5L  � �__s Q�  �x�]  5P�  Ru�]  �g�]  � i�7  5p�  �j�  u�7  �x�6  5��  �u�6  �x�6  5��  -u�6  �   m�W  O   ���  g�W  � g�W  � dO   h�W  	 i�7  X��  ��  g�7  ( w�6  X   �g�6  ( w�6  X   -g�6  (    rj�U    rO�    .5  �U  =�   �   ��   >�  �B  ?�  ��  EF�   �   �B   FF�  �C  GF�  �e  HF�  �8  IF�  ��  JF�  �

  X��   �   ��  Y��  ��
  Z��  ��   `Ŗ  �   ��  fז   �   ��  gז  ��  hז  ��  n�   �   ��	  o�  ��  p�  �H  v/�   �   �`  w/�  �w  x/�  �   y/�  �~  h�   �   �   �h�  ��  �h�  �  �h�  ��   �h�  ��  �h�  ��	  �h�  ��  �ȗ   �   �  �ȗ  �  �ȗ  ��  �ȗ  ��  ��   �   ��  ��  ��  ��  ��  ��  �m  �:�     �	  �:�  �2	  �:�  ��  �:�  �9  �:�  �[  ���     �J  ���  ��  ���  �7  ���  ��  ���     �I	  ���  �$	  ���  ��   ��   "  �N  ��  �p  ��   -  ��  ��  �:  ��  ��  ��  �d   ��  ��  �J�   8  �  �J�  ��  �J�  ��	  �v�   C  ��  �v�  �  ؕ�   N  ��  ٕ�  ��  ڕ�  ��  ە�  �+  �Ι   Y  ��  �Ι  ��   �Ι  �  ���   d  ��
  ���  ��  ���  �  �&�   o  �   �&�  �F  �&�  ��  �R�   z  ��  �R�  ��  �R�  �D  O~�   �  ��  P~�  �1  Q~�  ��  W��   �  �^  X��  ��  3ɚ   �  ��  4ɚ  ��   8�   �  ��  9�  �l	  =�  �  �N  >�  �^  ?�  �L  @�  �a  D@�  �  �B  E@�  ��	  F@�  �  G@�  �  H@�  �y  I@�  ��   ��   �  ��  !��  �  $�1  ��  �   �>  Y  �    9?   ^Y  �5 ,/ �V  x�      ��  (  �  �  �  E   �  �  o  �	  �  qW  !s   int   "�   �  #  .  <h   `  Ds   �  Wh   �  _z   �  es   t   ms   a  us     ~s   �  �s   3  �s   �  �s   H  �s   y  �s     �s   s  �s   T   �s   �  �s   F  �s   �  �s   �  �s     �s   V  �s   3   �  s  N:   �  V:   \	  2s   o  7s   �  <s   �  Cs   �  s   �  �  3   		pO qO 	!�  
std  �+  @�  %  0�=  
��  �b  
�3   Fe  
�s   �3  
�=  [  �-  �-   +  eq 
�<-  �-  }  �-  �-   lt 
��1  �-  �  �-  �-   ��  
eF  s   �  �-  �-  �   �K  
�9  �  �  �-   �(  

!  �-  �  �-  �  �-   1  
�A  �-     �-  �-  �   �5  
�'  �-  D  �-  �-  �   �3  
�A  �-  h  �-  �  +   +  
:  +  �  �-   6  �C  
 �P  6  �  �-   �B  
$6  �-  �  �-  �-   eof 
(�:  6  ?  
,N0  6  �-    _� �,   5�-  6�.  7/  �?  �%   K  \�  �+   �e  _�  �4  c,/  �J  d2/  ��  qY  _  J/   ��  so  z  J/  P/   W  y�  J/  s       �J  p  �B  �     %  �   �B  �  g/  �  P/    �e  y%  [V  �  �  �G  !�   <  x  �4  {1  �J  |=  �J  A-  `S  �F-  ~J  �  �J  �  �%  ��  �K  ��   I  ��  :!  �!/   %H  �D  _    �3  2�   �G  7�   t3  B�/  !�'  ��O  /  "V  ��N  �-  �  �  �/   "3  �o+  �-      �/   #�P  ��O    %  y/   #�M  ��P  8  >  y/   #�,  �-  Q  \  y/  �   "�+  ��R  �  s  y  y/   "3  �   �  �  �  y/  P/  P/   �/  !�B  y/  �  �  �  P/   #�O  �|6  �  �  y/  P/   $(  ��6  �    y/  P/   %�   �-  �      y/   &�1  o�*  �  3  y/  P/  �    %�A  $n%  �  \  b  m/   %�A  (�I  �  z  �  s/  �   %"A  ,�%  y/  �  �  m/   %�1  2E)  /  �  �  m/   %�/  6;&  /  �  �  m/   $�>  :�>  �  �  s/   %S  A:2  �    !  m/  �  �   $�#  K�(  5  J  m/  �  �  �   %9  S>$  �  b  r  m/  �  �   %-U  [�7  �-  �  �  m/  �   '�5  d�-  �  �  �  �   '	1  m�P  �  �  �  �   '�3  v\-  �  �  �  3    'nU  ��-  	  �  /  /   'nU  �nG  5	  �  ;  ;   'nU  ��   U	  �  �  �   'nU  �IP  u	  �  �  �   �J  �rR  s   �	  �  �   $�=  ��H  �	  �	  s/  �  �  �   $V  �)  �	  �	  s/   (�'  �D*  /  )�0  ��	  �	  s/   *�0  �
  
  s/  P/   �0  �)
  4
  s/  �/   �0  �D
  Y
  s/  �/  �  �   �0  �i
  �
  s/  �/  �  �  P/   �0  ��
  �
  s/  �  �  P/   �0  ��
  �
  s/  �  P/   �0  ��
  �
  s/  �  3   P/   )�0  "�
  	  s/  s    +�  *,Q  �/  "  -  s/  �/   +�  2�G  �/  F  Q  s/  �   +�  =�%  �/  j  u  s/  3    +S� f�&  /  �  �  s/   +S� q�>  ;  �  �  m/   ,end y<  /  �  �  s/   ,end �6;  ;  �  �  m/   +I ��$  S  
    s/   +I ��7  G  )  /  m/   +��  �lC  S  H  N  s/   +��  �CM  G  g  m  m/   +r ��R  �  �  �  m/   +�K  �r5  �  �  �  m/   +�3  �j=  �  �  �  m/   -�� �  �  �  s/  �  3    -�� ��F      s/  �   +I  v  �  (  .  m/   -�E  �|U  C  N  s/  �   -�1  -�  c  i  s/   +�� 5�?  �-  �  �  m/   +�:  D�6  #  �  �  m/  �   +�:  UW    �  �  s/  �   ,at k
/  #  �  �  m/  �   ,at ��7        s/  �   +�F  ��/  �/  /  :  s/  �/   +�F  �k:  �/  S  ^  s/  �   +�F  ��H  �/  w  �  s/  3    +@  DA:  �/  �  �  s/  �/   +@  U�1  �/  �  �  s/  �/  �  �   +@  )�D  �/  �  �  s/  �  �   +@  ��*  �/    !  s/  �   +@  �6  �/  :  J  s/  �  3    -�G  -aN  _  j  s/  3    .�3  �b*  �/  �  �  s/  �/   +�3  ^ 2  �/  �  �  s/  �/  �  �   +�3  �=  �/  �  �  s/  �  �   +�3  z�T  �/  �    s/  �   +�3  � @  �/  !  1  s/  �  3    -� ��E  F  [  s/  /  �  3    +� �\+  �/  t  �  s/  �  �/   +� �u>  �/  �  �  s/  �  �/  �  �   +� g|=  �/  �  �  s/  �  �  �   +� "�@  �/  �    s/  �  �   +� 9k<  �/  '  <  s/  �  �  3    +� K�'  /  U  e  s/  /  3    +bL  d�R  �/  ~  �  s/  �  �   +bL  t�2  /  �  �  s/  /   +bL  �L&  /  �  �  s/  /  /   +�%  �9F  �/  �  	  s/  �  �  �/   +�%  �|<  �/  "  A  s/  �  �  �/  �  �   +�%  ��T  �/  Z  t  s/  �  �  �  �   +�%  ��A  �/  �  �  s/  �  �  �   +�%  b>  �/  �  �  s/  �  �  �  3    +�%  3%  �/  �    s/  /  /  �/   +�%  'V7  �/    6  s/  /  /  �  �   +�%  <�+  �/  O  d  s/  /  /  �   +�%  Q'S  �/  }  �  s/  /  /  �  3    +�%  vj.  �/  �  �  s/  /  /  �  �   +�%  ��9  �/  �  �  s/  /  /  �  �   +�%  �C  �/    0  s/  /  /  /  /   +�%  �>/  �/  I  c  s/  /  /  ;  ;   %�?  ��&  �/  {  �  s/  �  �  �  3    %�1  �O  �/  �  �  s/  �  �  �  �   ,)  �z-  �  �  �  3   P/   /+E  �3J  �    �  3   P/   +�5  ��)  �  '  <  m/  �  �  �   -n	 @D  Q  \  s/  �/   +W�  �6  �  u  {  m/   +�A  %�A  �  �  �  m/   +��  ,Z5    �  �  m/   +�(  �;  �  �  �  m/  �  �  �   +�(  I�%  �       m/  �/  �   +�(  X�5  �  )  9  m/  �  �   +�(  �^   �  R  b  m/  3   �   +�(  v�S  �  {  �  m/  �/  �   +�(  	K  �  �  �  m/  �  �  �   +�(  �o?  �  �  �  m/  �  �   +�(  J5  �  �    m/  3   �   +NW  ��Q  �  $  4  m/  �/  �   +NW  /�I  �  M  b  m/  �  �  �   +NW  ��,  �  {  �  m/  �  �   +NW  ��;  �  �  �  m/  3   �   +�S  ��I  �  �  �  m/  �/  �   +�S  >T?  �  �    m/  �  �  �   +�S  05  �  $  4  m/  �  �   +�S  $S:  �  M  ]  m/  3   �   +�>  2hL  �  v  �  m/  �/  �   +�>  SUB  �  �  �  m/  �  �  �   +�>  Q�2  �  �  �  m/  �  �   +�>  _�K  �  �    m/  3   �   +�4  qT  �    /  m/  �/  �   +�4  j�K  �  H  ]  m/  �  �  �   +�4  ��5  �  v  �  m/  �  �   +�4  N.  �  �  �  m/  3   �   +U+  �)  �  �  �  m/  �  �   +��  �!1  s   �  �  m/  �/   +��  ��T  s     *  m/  �  �  �/   +��  ��O  s   C  b  m/  �  �  �/  �  �   +��  �;.  s   {  �  m/  �   +��  ��B  s   �  �  m/  �  �  �   +��  ��,  s   �  �  m/  �  �  �  �   �  0!T  3   1�E    1�F     2�&  2�7  �  �o  >�   �| Cs   3Q  b<   #  3�F c<  3�R  d<  33  e<  3�  f<  3�K  g<  3�@  h<   4all i<  ?5�� ��  :!  �!/   NF  ��/  �E  ��  p0  ��/  �%  ��/  6S  ��/  6�R  ��/  63  ��/  6�$  ��/  6�K  ��/  6�@  ��/  6�@  ��/  $�4  �Z  S  Y  �/   $�=  y)  m  s  �/   7�� �  �  �/  0  �   7�� �  �  �/  �  �   7�� �  �  �/  �   7N  �  �  �/  s    7�� �    �/  0   $�  �U    #  �/  0   %�&  �.  �-  ;  A  �/   $�F  &�;  U  e  �/  0  #   $�9  )�Q  y  �  �/  0  0   $WR  ,`2  �  �  �/  0  �/   $�S  /=  �  �  �/  �/  �/   8e  7,  �  �/  �/  �    �$  �/   6OD  �/  6gP  �/  6�F  $�/  2< 9id ��  �U  ��   6�I  �!/  $�  �<?  b  m  �/  �/   :id �|  �  �/  �/   ;id ��  �  �/   <4H  ��(  �  �  �/    �o  u�  �  �/   �o  ~�  �  �/  �/   *�o  ��    �/  �   �o  �  *  �/  �/  �  #   �o  �:  O  �/  �/  �/  #   5  �_  j  �/  s    .�  ��*  �/  �  �  �/  �/   .H�  ��N  �   �  �  �/   .U  �9  �-  �  �  �/  �/   .2  �t*  �-  �  �  �/  �/   =jP  �D       �/   >RD  �Q  �/  ?�o  7-   8   �/  �/   @�K  :�N  @�A  =�5  �K  @I  #  j   #   $�,  CH<  ~   �   �/  �/  �/  #   (  #  �     � >�  AW  3B!  B�4  B�$  Bq-  Bc=  Bo'  B�5   B�%  � B�8  �BX)  �B�%  �B�  �BaO  �BY=  � BP  �� B�C  ��BwS  �B�O  � B�?  �B�5  �� A
$ g{!  B)W  B�   B�U  B�A  B�8  B�P   BEH  �� A�4  ��!  BO   B�7  B(  B�Q  BG  �� A��  ��!  B�R   B�-  B�1  BlO  �� Cb4 p��!  )  D�3 � "  B�3  Bx0 BC5  E�3 ��"  '5 �0   � ��"  �U  �s   :!  �!/  7�3 �R"  g"  0  �"  s   0   $�4  ��2 {"  �"  0   &�=  �]- s   �"  0    F>. �!0  E�4 ��"  ?6 ��   �+ �%   �4 ��"  B0    G��"  B�0  5u�  K#  6�I  !/  6W�  �-  )u�  ,#  2#  H0   Ht�  ?#  H0  s     I\4 _0   �P  ��   J�4  p#  V#  Kdec p#  Jt-  p#  Khex p#  Jr'  p#  J< p#   Koct p#  @J� p#  �L[)  p#   L�%  "p#   L�  &p#   LdO  )p#   L\=  ,p#   L�P  /p#    L�C  3p#   @JzS  6p#  �J�O  9p#  JL�?  <p#  F�  J{!  J�7  N�$  k$  J(  Q�$  J�Q  V�$  JO  Y�$   F�9  iB!  Kapp l�$  �$  Kate o�$  J@� t�$  Kin w�$  Kout z�$  J�P  }�$   F�N  ��!  Kbeg �5%   %  Kcur �5%  Kend �5%  M�/ �+  Mi6 �+  Mk4 �V#  M�. �k$  M, �k$  M3 �0  M=4 ��"  M�1  o0  $M
. s   dM�- B0  hM*- 
  lNT3 m�0 &  &  0  �"  s    N8- �'3 (&  3&  0  �!   N/ �. G&  M&  0   .Q5 rH6 �0  e&  u&  0  s   �-   -f3 �, �&  �&  0   +n4 '�T  V#  �&  �&  �0   +n4 2�t  V#  �&  �&  0  V#   +s0 B?  V#  �&  �&  0  V#   +s0 S�(  V#  '   '  0  V#  V#   -q0 b�1 5'  @'  0  V#   +�/ m��  +  Y'  _'  �0   +�/ v2  +  x'  �'  0  +   +l6 ��K  +  �'  �'  �0   +l6 �6N  +  �'  �'  0  +   =d�  �c�  �-  �'  �-   +�= ��,   �'  (  0  �/   +-H  ��`    (  $(  �0   +*H  ��7  �/  =(  C(  �0   Or. d�- s   +�+ ��4 �0  l(  w(  0  s    +B6 ��0 �0  �(  �(  0  s    PS- W�!  �(  �(  0  s    b4 L�(  �(  0   7b4 �(  �(  0  N0   &�  <1 <0   )  0  N0    �!  A�0 �<)  BR1 B�1  B�1 B�2 B�3  AF2 �[)  B/ Bv/  B�4  <)  )  F0 �+  Q�+ �b/  Q}�  �]/  Q�. �]/  	Q�3 �b/  Q�. �b/  QJ- �b/  Q_5 �]/  Q�4 �]/   Qr6 �]/   Qf1 �]/   Q0 �]/   Q/, �b/   Q�1 �b/   QY2 �b/   QV, �[)   Q5 �b/   Qx, b/   Q�+ b/  Q�2 b/   Q�4 b/  Q�3 b/   Q�0 `)   min �n3 s   max ��, s   (T4 �2 s   (/5 ��. s   (�2 �2 s   (�1 M. s   (]2 �3 s   (�4 s1 s    �>  b  R�*  �{!  6+  {!  {!   R	W  �w1  P+  }1  {!   {!  R*  �{!  o+  {!  {!   2z o+  St4 _�/ �    T$   �|-  �  $,�  -  K  :<-  �e  =�  � ?�  "  @�  �4  A,/  �J  B2/  �A  O,  	,  8/   �A  Q,  $,  8/  >/   �A  V4,  ?,  8/  s    .�
 Y51  �+  W,  b,  D/  �+   .�
 ]�R  �+  z,  �,  D/  �+   .� c?  �+  �,  �,  8/  �+  �   N_ m.   �,  �,  8/  �+  �+   .�3  q89  �+  �,  �,  D/   N.E  ��3  -  -  8/  �+  2/   N�(  ��(  '-  2-  8/  �+   U_Tp 3    �+  2ZD  28E  VU  A!/  e-  �0  s    W9+  N!/  �0  s     �� �� �� T2*  7�-  X8   Y+  Y[  �  [  +  Y�  �  8�.  �{  �   ]�  �  \�   �  �D  !�  �3  "�  U>  #�  &�  $�  �  %�  �*  &�   ڡ  '3   $�U  (3   %TL  )3   &�I  *3   'Q  +3   (�C  ,3   )�J  -3   *1  .�  ,o(  /3   0�U  03   1PL  13   2�I  23   3Q  33   4�C  43   5�J  53   6 R)%  K�  /  s   �   ZGT  P/  �-  �   s   Y3   Y�  �+  Y<-  <-    Y�    s   �-  �    �  �  Y�  Y  Y�  [,   �/  \ �  �  �/  �/  �    Y�   �   (  Y�   �   �/  �   �  [�/  �/  \ [0  0  \ 
0  �/  Y�   �    "  '0  ]<0  �!  <0  s    Y�!  �"  �"  Y)  ^s   _0  _ e0  `�5  T0  [�"  0  a�   �!  Y�"  )  Y%   Y�  !/  bK-  �0  cXF  A�0  c\;  As   de�T  C!/    b+  �0  f__a �{!  f__b �{!   be-  1  cXF  N�0  c\;  Ns    g�"  !1  +1  hh  +1   B0  gB"  >1  l1  hh  l1  iJ4 ��"  i;5 �s   i�1 �0   0  j�*  YP+  Y{!  b6+  �1  f__a ��1  f__b �{!   }1  bU+  �1  f__a �{!  f__b �{!   g�"  �1  �1  hh  l1  dk/t  �s     g�(   �1  2  hh  2   0  l�1  c/ p{   �(2  q2  m�1  = n1  �   ON2  m!1  _  n1  �   Ok2  m!1  �  o� pC(  �   ��2  q�   r#- h!/  �Es�0  ���  it1  u�0  �E�s�0  ���  Vt�0  u�0  �E�v��  w�0  �      x�%   1   �
3  p3  yh  2  � zJ4 m�"  �z;5 ms   �n01      nf3  m_1  � uS1  �uG1  �u>1  P { �>   xM&  P �  ��3  5  yh  2  � zO4 rs   �z�3 r�-  �|��  �4  }<2 us   � }3 vB0  q n1  �    }�3  m!1  �  ~� ;   4  __i �s     ~�!`   �4  �5  ��1  �!��  �f4  t�1  m�1  ' s�0  �!�  �t�0  m�0  L   {�!�>  {�!�>  {�!y+  {�!�>   ��1  @! �  ��4  m�1  ` m�1  � ��0  @!   �m�0  ` m�0  �   {� �>  {!�>  {�!y+   {�!?  {�!?   	5  Yt+  �&   "f   �'5  �5  yh  2  � �__e ��!  �|8�  m5  __p �0  � {E"�>  {M"�>   {]"?  {f"?   x3&  p"]   ��5  ^6  yh  2  � qy"N   __p �0   ��1  �"P�  �:6  m�1   vP�  ��1  ��0  �"P�  �m1  = m�0  R s�0  �"P�  Vm�0  = m�0  R vP�  w�0  t      q�"   }4 �0  � {�"+?     g�(   l6  6  hh  2  h#  ]/   l^6  �1 �"R   ��6  �6  ul6  � {�"5  {�"�5  {#�>  o"# l^6  }5 0#   ��6  �6  ul6  � {>#6  �K#+?   �U  =7   �   ��   >7  �B  ?7  ��  E37   �   �B   F37  �C  G37  �e  H37  �8  I37  ��  J37  �

  X�7   �   ��  Y�7  ��
  Z�7  ��   `�7  �   ��  f�7   �   ��  g�7  ��  h�7  ��  n�7   �   ��	  o�7  ��  p�7  �H  v8   �   �`  w8  �w  x8  �   y8  �~  U8   �   �   �U8  ��  �U8  �  �U8  ��   �U8  ��  �U8  ��	  �U8  ��  ��8   �   �  ��8  �  ��8  ��  ��8  ��  ��8   �   ��  ��8  ��  ��8  ��  ��8  �m  �'9     �	  �'9  �2	  �'9  ��  �'9  �9  �'9  �[  �m9     �J  �m9  ��  �m9  �7  �m9  ��  ��9     �I	  ��9  �$	  ��9  ��   ��9   "  �N  ��9  �p  ��9   -  ��  ��9  �:  ��9  ��  ��9  �d   ��9  ��  �7:   8  �  �7:  ��  �7:  ��	  �c:   C  ��  �c:  �  ؂:   N  ��  ق:  ��  ڂ:  ��  ۂ:  �+  �:   Y  ��  �:  ��   �:  �  ��:   d  ��
  ��:  ��  ��:  �  �;   o  �   �;  �F  �;  ��  �?;   z  ��  �?;  ��  �?;  �D  Ok;   �  ��  Pk;  �1  Qk;  ��  W�;   �  �^  X�;  ��  3�;   �  ��  4�;  ��   8�;   �  ��  9�;  �l	  =�;  �  �N  >�;  �^  ?�;  �L  @�;  �a  D-<  �  �B  E-<  ��	  F-<  �  G-<  �  H-<  �y  I-<  ��   �<   �  ��  !�<  �b#  <, �		�u#  �+ �		��#  �/ �		��#  �. �		��#  , �		��#  - �		��#  �. �		��#  k2 �		��#  �0 �		��#  �- �		��#  ,0 �		�$  e5 �		�$  �, �		�"$  �4 |		�1$  �2 x		�@$  �/ t		�N$  0 p		�\$  �, l		�x$  Z0 h		��$  �+ d		��$  �4 `		��$  y. \		��$  )4 X		��$  �0 T		��$  a, P		��$  �- L		��$  �4 H		�%  &1 D		�'%  4 @		�:%  �5 <		�H%  �5 8		�#  H�/ �E�#  J�- hD/�  ��  �  �>  �   ��  �  �>  �   ��  /�  ��  �  �>  �   �e  �Ӫ  ?  �   �>  Y  ?  �   �  +?  �   S�  �1  �    �/   �a  �6 �7 �V  H�      P�  (  _� �7   �  �  8k  �{  k   ]�  k  \�   k  �D  !k  �3  "k  U>  #k  &�  $k  �  %k  �*  &k   ڡ  'q  $�U  (q  %TL  )q  &�I  *q  'Q  +q  (�C  ,q  )�J  -q  *1  .k  ,o(  /q  0�U  0q  1PL  1q  2�I  2q  3Q  3q  4�C  4q  5�J  5q  6 q  �  std  n  5>   6n  7�  @R!  	%  0�=  �n  �b  �q  Fe  �  
�3  �=  �  e%  k%   �  eq �<-  q%    k%  k%   lt ��1  q%  !  k%  k%   ��  eF  �  E  x%  x%  n   �K  �9  n  _  x%   �(  
!  x%  �  x%  n  k%   1  �A  ~%  �  ~%  x%  n   �5  �'  ~%  �  ~%  x%  n   �3  �A  ~%  �  ~%  n  �   +  :  �  	  �%   �  �C   �P  �  (  k%   �B  $6  q%  G  �%  �%   eof (�:  �  ?  ,N0  �  �%    _� 	�7   �?  	�%   K  
\  }!   �e  
_n  �4  
c�%  �J  
d�%  ��  
q�  �  �%   ��  
s�  �  �%  �%   W  
y�  �%  �    �  �J  pz  �B  R  �   %  k   �B  A  �%  k  �%    �e  y�  [V  k  R  �G  !   <  x�  �4  {�  �J  |�  �J  #  `S  �2%  ~J  �z  �J  �  �%  �  �K  �R   I  �R  :!  ��%   %H  ��  �   �3  2k  �G  7�  t3  B�%  �'  ��O  �%  V  ��N  q%  [  a  �%   3  �o+  q%  x  ~  �%   �P  ��O  �  �  �%   �M  ��P  �  �  �%   �,  �-  �  �  �%  R   �+  ��R  k  �  �  �%   3  �   k      �%  �%  �%   �/  !�B  �%  6  R  R  �%   �O  �|6  I  T  �%  �%    (  ��6  h  s  �%  �%   !�   �-  k  �  �  �%   "�1  o�*  k  �  �%  �%  R    !�A  $n%  k  �  �  �%   !�A  (�I  k  �  �  �%  k   !"A  ,�%  �%      �%   !�1  2E)  �  -  3  �%   !�/  6;&  �  K  Q  �%    �>  :�>  e  k  �%   !S  A:2  R  �  �  �%  R  �    �#  K�(  �  �  �%  R  R  �   !9  S>$  R  �  �  �%  R  R   !-U  [�7  q%  �    �%  �   #�5  d�-  '  k  �  R   #	1  m�P  G  k  �  R   #�3  v\-  g  k  R  q   #nU  ��-  �  k  �  �   #nU  �nG  �  k  �  �   #nU  ��   �  k  k  k   #nU  �IP  �  k  �  �   �J  �rR  �  	  R  R    �=  ��H  	  /	  �%  R  R  R    V  �)  C	  I	  �%   $�'  �D*  �%  %�0  �j	  p	  �%   &�0  ��	  �	  �%  �%   �0  ��	  �	  �%  �%   �0  ��	  �	  �%  �%  R  R   �0  ��	  �	  �%  �%  R  R  �%   �0  �
  
  �%  �  R  �%   �0  �*
  :
  �%  �  �%   �0  �J
  _
  �%  R  q  �%   %�0  "p
  {
  �%  �   '�  *,Q  �%  �
  �
  �%  �%   '�  2�G  �%  �
  �
  �%  �   '�  =�%  �%  �
  �
  �%  q   'S� f�&  �       �%   'S� q�>  �    %  �%   (end y<  �  >  D  �%   (end �6;  �  ]  c  �%   'I ��$  �  |  �  �%   'I ��7  �  �  �  �%   '��  �lC  �  �  �  �%   '��  �CM  �  �  �  �%   'r ��R  R  �  �  �%   '�K  �r5  R      �%   '�3  �j=  R  6  <  �%   )�� �  Q  a  �%  R  q   )�� ��F  v  �  �%  R   'I  v  R  �  �  �%   )�E  �|U  �  �  �%  R   )�1  -�  �  �  �%   '�� 5�?  q%  �  �  �%   '�:  D�6  �      �%  R   '�:  UW  �  7  B  �%  R   (at k
/  �  Z  e  �%  R   (at ��7  �  }  �  �%  R   '�F  ��/  �%  �  �  �%  �%   '�F  �k:  �%  �  �  �%  �   '�F  ��H  �%  �  �  �%  q   '@  DA:  �%      �%  �%   '@  U�1  �%  1  F  �%  �%  R  R   '@  )�D  �%  _  o  �%  �  R   '@  ��*  �%  �  �  �%  �   '@  �6  �%  �  �  �%  R  q   )�G  -aN  �  �  �%  q   *�3  �b*  �%  �  �  �%  �%   '�3  ^ 2  �%    -  �%  �%  R  R   '�3  �=  �%  F  V  �%  �  R   '�3  z�T  �%  o  z  �%  �   '�3  � @  �%  �  �  �%  R  q   )� ��E  �  �  �%  �  R  q   '� �\+  �%  �  �  �%  R  �%   '� �u>  �%    )  �%  R  �%  R  R   '� g|=  �%  B  W  �%  R  �  R   '� "�@  �%  p  �  �%  R  �   '� 9k<  �%  �  �  �%  R  R  q   '� K�'  �  �  �  �%  �  q   'bL  d�R  �%  �     �%  R  R   'bL  t�2  �    $  �%  �   'bL  �L&  �  =  M  �%  �  �   '�%  �9F  �%  f  {  �%  R  R  �%   '�%  �|<  �%  �  �  �%  R  R  �%  R  R   '�%  ��T  �%  �  �  �%  R  R  �  R   '�%  ��A  �%  �    �%  R  R  �   '�%  b>  �%  -  G  �%  R  R  R  q   '�%  3%  �%  `  u  �%  �  �  �%   '�%  'V7  �%  �  �  �%  �  �  �  R   '�%  <�+  �%  �  �  �%  �  �  �   '�%  Q'S  �%  �  	  �%  �  �  R  q   '�%  vj.  �%  "  <  �%  �  �  k  k   '�%  ��9  �%  U  o  �%  �  �  �  �   '�%  �C  �%  �  �  �%  �  �  �  �   '�%  �>/  �%  �  �  �%  �  �  �  �   !�?  ��&  �%  �    �%  R  R  R  q   !�1  �O  �%    9  �%  R  R  �  R   ,)  �z-  k  ]  R  q  �%   ++E  �3J  k  �  R  q  �%   '�5  ��)  R  �  �  �%  k  R  R   )n	 @D  �  �  �%  �%   'W�  �6  �  �  �  �%   '�A  %�A  �      �%   '��  ,Z5  }  %  +  �%   '�(  �;  R  D  Y  �%  �  R  R   '�(  I�%  R  r  �  �%  �%  R   '�(  X�5  R  �  �  �%  �  R   '�(  �^   R  �  �  �%  q  R   '�(  v�S  R  �  �  �%  �%  R   '�(  	K  R    +  �%  �  R  R   '�(  �o?  R  D  T  �%  �  R   '�(  J5  R  m  }  �%  q  R   'NW  ��Q  R  �  �  �%  �%  R   'NW  /�I  R  �  �  �%  �  R  R   'NW  ��,  R  �  �  �%  �  R   'NW  ��;  R    &  �%  q  R   '�S  ��I  R  ?  O  �%  �%  R   '�S  >T?  R  h  }  �%  �  R  R   '�S  05  R  �  �  �%  �  R   '�S  $S:  R  �  �  �%  q  R   '�>  2hL  R  �  �  �%  �%  R   '�>  SUB  R    &  �%  �  R  R   '�>  Q�2  R  ?  O  �%  �  R   '�>  _�K  R  h  x  �%  q  R   '�4  qT  R  �  �  �%  �%  R   '�4  j�K  R  �  �  �%  �  R  R   '�4  ��5  R  �  �  �%  �  R   '�4  N.  R    !  �%  q  R   'U+  �)  	  :  J  �%  R  R   '��  �!1  �  c  n  �%  �%   '��  ��T  �  �  �  �%  R  R  �%   '��  ��O  �  �  �  �%  R  R  �%  R  R   '��  �;.  �  �  �  �%  �   '��  ��B  �    &  �%  R  R  �   '��  ��,  �  ?  Y  �%  R  R  �  R     ,!T  q  -�E  �  -�F  �   .�&  .�7  	  � >	  /W  3#  0�4  0�$  0q-  0c=  0o'  0�5   0�%  � 0�8  �0X)  �0�%  �0�  �0aO  �0Y=  � 0P  �� 0�C  ��0wS  �0�O  � 0�?  �0�5  �� /
$ g\  0)W  0�   0�U  0�A  0�8  0�P   0EH  �� /�4  ��  0O   0�7  0(  0�Q  0G  �� 1b4 0  'n4 '�T  �  �  �  �'   �P  ��  2�4  �  �  3dec �  2t-  �  3hex �  2r'  �  2< �   3oct �  @2� �  �4[)  �   4�%  "�   4�  &�   4dO  )�   4\=  ,�   4�P  /�    4�C  3�   @2zS  6�  �2�O  9�  J4�?  <�  5�  J\  2(  Q�  �  2�Q  V�  2O  Y�   5�9  i#  3in w    3out z   6;v  ��  7��  09�   0�  0�  0˭  0�  0^�  0j  0L�  $0ڭ  0<�  "03�  $ Ў  �  r  �  86�  �k  &  k  q    �  <&  =&  >"&  @�&  A�&  B�&  C�&  D'  E-'  FM'  Gb'  Hw'  6�  H�  9�k  KU  0Q   0� 0ʄ  0ih  0~  :Sv  Lq  �O  L�'    �  N~  U  ��  Y�  ;Fv  ^��  U  q  q  q    ד  ��  ��  �y  � �k  �4  ��%  ,{�  k   <*  K�    �  �   <ͳ  �Y(  &  =_Tp 7   Y(  Y(   +��  [Ki  q%  I  �  n  [)   �  n  >�  �   �/  ,!T  q    <)%  Kk  �  �  �   ?int �  q  @GT  P�  >   �  �  �  �  o  �	  �  qW  !�    "�  �  #  .  <�  `  D�  �  W�  �  _�  �  e�  t   m�  a  u�    ~�  �  ��  3  ��  �  ��  H  ��  y  ��    ��  s  ��  T   Ȉ  �  Ј  F  ׈  �  ��  �  �    �  V  �  �  s  N�  �  V�  \	  2�  o  7�  �  <�  �  C�  �  �  I!  ABpO qO !J!  C$   E=%  	�  $,n  -y  K  :#  �e  =n  � ?k  "  @�  �4  A�%  �J  B�%  �A  O�!  �!  �%   �A  Q�!  �!  �%  �%   �A  V"  "  �%  �   *�
 Y51  �!  )"  4"  �%  �!   *�
 ]�R  �!  L"  W"  �%  �!   *� c?  �!  o"  "  �%  �!  C!   D_ m.   �"  �"  �%  �!  �!   *�3  q89  �!  �"  �"  �%   D.E  ��3  �"  �"  �%  �!  �%   D�(  ��(  �"  #  �%  �!   =_Tp q   }!  6ZD  �2%  EF�  �k   5��  ��  5�4  ��  5� ��  %��  �f#  l#  �'   F��  �}#  �#  �'  �'   '*  ��}  ;#  �#  �#  �'   'Ư  �?s  H#  �#  �#  �'   '�F  �Ϭ  �'  �#  �#  �'   '�F  ��  #  �#  	$  �'  �   'a�  �
�  �'  "$  ($  �'   'a�   ��  #  A$  L$  �'  �   '�:  ,�  ;#  e$  p$  �'  .#   '�F  		n  �'  �$  �$  �'  .#   '(*  ��  #  �$  �$  �'  .#   ' I  h�  �'  �$  �$  �'  .#   '�O  7k  #  �$   %  �'  .#   'WC  ]�  �'  %  %  �'   ,{�  k  ,�  	   .8E  #   �� �� �� C2*  7e%  G8�   H�  H�  �  �  �  H	  Hq  H�  }!  H#  #  �  H    �   �    �  	    H  H�  H	  I7   �%  J Y  7   H�  �l  %   j�  #%   Ktm ,,�&  ,g  .�   �  /�  �  0�  ��  1�  ��  2�  ��  3�  ��  4�  �  5�  d�  6�   ��  7%   $~�  8�  ( @\�  >&  <ѯ  HD%  �&  &  &   <��  M&  �&  �&   "&  <�  C&  '  '   &  <#�  ak  "'  "'   ('  "&  <�� fk  B'  B'   H'  &  <��  W�&  b'  B'   <[v  \�&  w'  B'   <��  R,   �'  k  ,   �  "'   Iq  �'  L�    #  H�'  k  7%  H#  M�  �'  �'  Nh  �'   �%  M�  �'  �'  Nh  �'   �  M�  (  (  Nh  (   �'  O�  A(  P__a K�  P__b K�   M�  O(  Y(  Nh  �'   H&  O  �(  =_Tp 7   P__a (  P__b (   Y(  Y(  M�  �(  �(  Nh  �'  Q%  DR   R�  =P#�   �V)  S$  =V)  � T�6 =k  � S!�  >q  �U��  V��  @�  V�6 O�  W (  �#   O6)  X5(  Y*(  3  Z (  �#   TY5(  Q [*(     &  HI  \&  �#�   �F*  T�  [�  g T��  [n  � S)�  \F*  �U��  ]__n ^N  � V�~  _N  ]__i `n  
 ^�7 aq%  @ _A(  �# �  ^+*  `O(  �a�'  �#�  �`�'  �a�'  �#0�  -`�'  �   b�#)   ]__j fn  �    [)  cU  =W*   �  c�   >W*  cB  ?W*  c�  E�*      cB   F�*  cC  G�*  ce  H�*  c8  I�*  c�  J�*  c

  X�*      c�  Y�*  c�
  Z�*  d�   `�*     c�  f+   )   c�  g+  c�  h+  c�  n0+   4   c�	  o0+  c�  p0+  cH  vY+   ?   c`  wY+  cw  xY+  c   yY+  c~  �+   J   c   ��+  c�  ��+  c  ��+  c�   ��+  c�  ��+  c�	  ��+  c�  ��+   U   c  ��+  c  ��+  c�  ��+  c�  �,   `   c�  �,  c�  �,  c�  �,  cm  �Q,   k   c	  �Q,  c2	  �Q,  c�  �Q,  c9  �Q,  c[  ��,   v   cJ  ��,  c�  ��,  c7  ��,  c�  ��,   �   cI	  ��,  c$	  ��,  c�   ��,   �   cN  ��,  cp  �-   �   c�  �-  c:  �-  c�  �-  cd   �-  c�  �N-   �   c  �N-  c�  �N-  c�	  �w-   �   c�  �w-  c  ؔ-   �   c�  ٔ-  c�  ڔ-  c�  ۔-  c+  ��-   �   c�  ��-  c�   ��-  c  ��-   �   c�
  ��-  c�  ��-  c  �.   �   c   �.  cF  �.  c�  �D.   �   c�  �D.  c�  �D.  cD  Om.   �   c�  Pm.  c1  Qm.  c�  W�.   !  c^  X�.  c�  3�.   !  c�  4�.  c�   8�.   !  c�  9�.  cl	  =�.  "!  cN  >�.  c^  ?�.  cL  @�.  ca  D"/  -!  cB  E"/  c�	  F"/  c  G"/  c  H"/  cy  I"/  c�   o/   8!  c�  !o/  e�  7�7 lDe�  6�6 pDI�  �/  L�    fX  �7 �Deq  2�6 5
	e�  4�6 tD t]   �g  : += �V  ��      ��  (  _� �7   �  �  8k  �{  k   ]�  k  \�   k  �D  !k  �3  "k  U>  #k  &�  $k  �  %k  �*  &k   ڡ  'q  $�U  (q  %TL  )q  &�I  *q  'Q  +q  (�C  ,q  )�J  -q  *1  .k  ,o(  /q  0�U  0q  1PL  1q  2�I  2q  3Q  3q  4�C  4q  5�J  5q  6 q  �  std ' f#  5>   6f#  7�#  R�#  U�#  [�#  \�#  	v�%  	w�%  	{&  	�!&  	�=&  	�R&  	�g&  	��&  	��&  	��&  	��&  	�'  	�D'  	�d'  	��'  	��'  	��'  	��'  	��'  	��'  
@(  	M8 \a  
^ȹ    %  0�=  �0  �b  �q  Fe  �#  �3  �=  �  &.  ,.   t  eq �<-  2.  �  ,.  ,.   lt ��1  2.  �  ,.  ,.   ��  eF  �#    9.  9.  0   �K  �9  0  !  9.   �(  
!  9.  E  9.  0  ,.   1  �A  ?.  i  ?.  9.  0   �5  �'  ?.  �  ?.  9.  0   �3  �A  ?.  �  ?.  0  t   +  :  t  �  E.     �C   �P    �  ,.   �B  $6  2.  	  E.  E.   eof (�:    ?  ,N0    E.    _� �7   �?  �%   K  \�  G(   �e  _0  �4  cK.  �J  dQ.  ��  q�  �  i.   ��  s�  �  i.  o.   W  y�  i.  �#    F  �J  pT  	�B  ,  F   %  k   �B      �.  k  o.   �B     �.  �#    �e  yY  [V  E  ,  �G  !�   <  xF  �4  {e  �J  |q  �J  �)  `S  ��+  ~J  �T  �J  �Y  �%  ��  �K  �,   I  �,  :!  ��.   %H  ��  �   �3  2E  �G  7�#  t3  B�.   �'  ��O  �.  !V  ��N  2.  5  ;  �.   !3  �o+  2.  R  X  �.   "�P  ��O  k  q  �.   "�M  ��P  �  �  �.   "�,  �-  �  �  �.  ,   !�+  ��R  k  �  �  �.   !3  �   k  �  �  �.  o.  o.   �/  !�B  �.    ,  ,  o.   "�O  �|6  #  .  �.  o.   #(  ��6  B  M  �.  o.   $�   �-  k  e  k  �.   %�1  o�*  k    �.  o.  ,    $�A  $n%  k  �  �  �.   $�A  (�I  k  �  �  �.  k   $"A  ,�%  �.  �  �  �.   $�1  2E)  {      �.   $�/  6;&  {  %  +  �.   #�>  :�>  ?  E  �.   $S  A:2  ,  ]  m  �.  ,  �#   #�#  K�(  �  �  �.  ,  ,  �#   $9  S>$  ,  �  �  �.  ,  ,   $-U  [�7  2.  �  �  �.  �#   &�5  d�-  	  k  �#  ,   &	1  m�P  !	  k  �#  ,   &�3  v\-  A	  k  ,  q   &nU  ��-  a	  k  {  {   &nU  �nG  �	  k  �  �   &nU  ��   �	  k  k  k   &nU  �IP  �	  k  �#  �#   �J  �rR  �#  �	  ,  ,   #�=  ��H  �	  	
  �.  ,  ,  ,   #V  �)  
  #
  �.   '�'  �D*  �.  (�0  �D
  J
  �.   )�0  �Z
  e
  �.  o.   �0  �u
  �
  �.  �.   �0  ��
  �
  �.  �.  ,  ,   �0  ��
  �
  �.  �.  ,  ,  o.   �0  ��
  �
  �.  �#  ,  o.   �0  �    �.  �#  o.   �0  �$  9  �.  ,  q  o.   (�0  "J  U  �.  �#   *�  *,Q  �.  n  y  �.  �.   *�  2�G  �.  �  �  �.  �#   *�  =�%  �.  �  �  �.  q   *S� f�&  {  �  �  �.   *S� q�>  �  �  �  �.   +end y<  {      �.   +end �6;  �  7  =  �.   *I ��$  �  V  \  �.   *I ��7  �  u  {  �.   *��  �lC  �  �  �  �.   *��  �CM  �  �  �  �.   *r ��R  ,  �  �  �.   *�K  �r5  ,  �  �  �.   *�3  �j=  ,      �.   ,�� �  +  ;  �.  ,  q   ,�� ��F  P  [  �.  ,   *I  v  ,  t  z  �.   ,�E  �|U  �  �  �.  ,   ,�1  -�  �  �  �.   *�� 5�?  2.  �  �  �.   *�:  D�6  o  �  �  �.  ,   *�:  UW  c      �.  ,   +at k
/  o  4  ?  �.  ,   +at ��7  c  W  b  �.  ,   *�F  ��/  �.  {  �  �.  �.   *�F  �k:  �.  �  �  �.  �#   *�F  ��H  �.  �  �  �.  q   *@  DA:  �.  �  �  �.  �.   *@  U�1  �.       �.  �.  ,  ,   *@  )�D  �.  9  I  �.  �#  ,   *@  ��*  �.  b  m  �.  �#   *@  �6  �.  �  �  �.  ,  q   ,�G  -aN  �  �  �.  q   -�3  �b*  �.  �  �  �.  �.   *�3  ^ 2  �.  �    �.  �.  ,  ,   *�3  �=  �.     0  �.  �#  ,   *�3  z�T  �.  I  T  �.  �#   *�3  � @  �.  m  }  �.  ,  q   ,� ��E  �  �  �.  {  ,  q   *� �\+  �.  �  �  �.  ,  �.   *� �u>  �.  �    �.  ,  �.  ,  ,   *� g|=  �.    1  �.  ,  �#  ,   *� "�@  �.  J  Z  �.  ,  �#   *� 9k<  �.  s  �  �.  ,  ,  q   *� K�'  {  �  �  �.  {  q   *bL  d�R  �.  �  �  �.  ,  ,   *bL  t�2  {  �  �  �.  {   *bL  �L&  {    '  �.  {  {   *�%  �9F  �.  @  U  �.  ,  ,  �.   *�%  �|<  �.  n  �  �.  ,  ,  �.  ,  ,   *�%  ��T  �.  �  �  �.  ,  ,  �#  ,   *�%  ��A  �.  �  �  �.  ,  ,  �#   *�%  b>  �.    !  �.  ,  ,  ,  q   *�%  3%  �.  :  O  �.  {  {  �.   *�%  'V7  �.  h  �  �.  {  {  �#  ,   *�%  <�+  �.  �  �  �.  {  {  �#   *�%  Q'S  �.  �  �  �.  {  {  ,  q   *�%  vj.  �.  �    �.  {  {  k  k   *�%  ��9  �.  /  I  �.  {  {  �#  �#   *�%  �C  �.  b  |  �.  {  {  {  {   *�%  �>/  �.  �  �  �.  {  {  �  �   $�?  ��&  �.  �  �  �.  ,  ,  ,  q   $�1  �O  �.  �    �.  ,  ,  �#  ,   ,)  �z-  k  7  ,  q  o.   .+E  �3J  k  Z  ,  q  o.   *�5  ��)  ,  s  �  �.  k  ,  ,   ,n	 @D  �  �  �.  �.   *W�  �6  �#  �  �  �.   *�A  %�A  �#  �  �  �.   *��  ,Z5  W  �    �.   *�(  �;  ,    3  �.  �#  ,  ,   *�(  I�%  ,  L  \  �.  �.  ,   *�(  X�5  ,  u  �  �.  �#  ,   *�(  �^   ,  �  �  �.  q  ,   *�(  v�S  ,  �  �  �.  �.  ,   *�(  	K  ,  �    �.  �#  ,  ,   *�(  �o?  ,    .  �.  �#  ,   *�(  J5  ,  G  W  �.  q  ,   *NW  ��Q  ,  p  �  �.  �.  ,   *NW  /�I  ,  �  �  �.  �#  ,  ,   *NW  ��,  ,  �  �  �.  �#  ,   *NW  ��;  ,  �     �.  q  ,   *�S  ��I  ,    )  �.  �.  ,   *�S  >T?  ,  B  W  �.  �#  ,  ,   *�S  05  ,  p  �  �.  �#  ,   *�S  $S:  ,  �  �  �.  q  ,   *�>  2hL  ,  �  �  �.  �.  ,   *�>  SUB  ,  �     �.  �#  ,  ,   *�>  Q�2  ,    )  �.  �#  ,   *�>  _�K  ,  B  R  �.  q  ,   *�4  qT  ,  k  {  �.  �.  ,   *�4  j�K  ,  �  �  �.  �#  ,  ,   *�4  ��5  ,  �  �  �.  �#  ,   *�4  N.  ,  �  �  �.  q  ,   *U+  �)  �    $  �.  ,  ,   *��  �!1  �#  =  H  �.  �.   *��  ��T  �#  a  v  �.  ,  ,  �.   *��  ��O  �#  �  �  �.  ,  ,  �.  ,  ,   *��  �;.  �#  �  �  �.  �#   *��  ��B  �#  �     �.  ,  ,  �#   *��  ��,  �#    3  �.  ,  ,  �#  ,   �  /!T  q  0�E  h  0�F  F   1�&  1�7  �  �o  >�"  20  �;  �| C�#  3Q  b�     3�F c�  3�R  d�  33  e�  3�  f�  3�K  g�  3�@  h�   4all i�  ?5�� �N  :!  ��.   NF  �/  �E  �0  p0  �/  �%  ��'  6S  �/  6�R  �/  63  �/  6�$  �/  6�K  �/  6�@  �/  6�@  �/  #�4  �Z  �  �  �.   #�=  y)  �  �  �.   �� �  �  �.  2/  0   �� �    �.  �#  0   ��   *  �.  0   N  :  E  �.  �#   �� U  `  �.  2/   #�  �U  t    �.  2/   $�&  �.  2.  �  �  �.   #�F  &�;  �  �  �.  8/     #�9  )�Q  �  �  �.  8/  '/   #WR  ,`2  �  	  �.  8/  �.   #�S  /=    -  �.  �.  /   7e  7,  =  �.  /  0    �$  �.   6OD  �.  6gP  �.  6�F  $�.  8< R  
   9< B1   :!  X�.  8 � #  :C8 �h1  C ;�A  �=9 << r�  �  m1  0   =< �  �    m1  �#   >��  z�r  )  s1  �#   #   ?��  ~�   #  D  s1   >�h  �ܧ  [  s1   ?�< ��;  #  {   #  �#   @�m  �~�   #  @��  ܧ�  �#  #�4  �l; �  �  /   #�=  ��8 �  �  /   < ��  �  m1  y1   %�  �= 1  �  m1  y1    Aid ��   �U  �0   6�I  ��.  #�  �<?  D   O   �.  �.   Bid �^   i   �.  �.   Cid �y      �.   D4H  ��(  0  �   �.    �o  u�   �   �.   �o  ~�   �   �.  �.   )�o  ��   �   �.  �#   �o  ��   !  �.  �.  �#     �o  �!  1!  �.  �.  �.     5  �A!  L!  �.  �#   -�  ��*  �.  d!  o!  �.  �.   -H�  ��N  �"  �!  �!  �.   -U  �9  2.  �!  �!  �.  �.   -2  �t*  2.  �!  �!  �.  �.   ?jP  �D  c  �!  �.   ERD  �Q  �.  F�o  7"  "  �.  �.   G�K  :�N  G�A  =�5  �K  @I    L"     #�,  CH<  `"  u"  �.  �.  �.     
     �   c  � >�  <I/  =>/  >T/  @�/  A�/  B	0  C$0  D?0  E_0  F0  G�0  H�0  ד  � #  ��  �;  � �k  �4  �K.  /{�  k   W�  1R1  H}�  �	�-  O#  /!T  q  �.  �.   0  I�8 R#< �#    J)%  Kk  �#  �#  �#   Kint �#  q  LGT  P�#  >   J��  E�#  �#  �#  �#   J��  Uk  �#  �#   J��  Ok  �#  k  �#   J��  F,   $  k  �#  ,    �  $  �  �  o  �	  �  qW  !�#    "O$  �  #  Ms  N$  �  V$  .  <9$  `  D�#  �  W9$  �  _D$  �  e�#  t   m�#  a  u�#    ~�#  �  ��#  3  ��#  �  ��#  H  ��#  y  ��#    ��#  s  ��#  T   Ȁ#  �  Ѐ#  F  ׀#  �  ��#  �  �#    �#  V  �#  �  \	  2�#  o  7�#  �  <�#  �  C�#  �  �#  N*  �%  �  �#   Orem �#   +   �%  N#@  �%  �  $%    Orem %%    A  &�%  J� ��#  &  &    &  PJ�  >6&  6&  �#   �� J�  H�#  R&  �#   J�  I%   g&  �#   J�  �]$  �&  �&  �&  ,   ,   �&   �&  Q�&  R�#  �&  �&  �&   Sdiv �%  �&  �#  �#   J    �k  �&  �#   H�   �%  �&  %   %    H�  .�#  '  �#  ,    H�  \,   7'  7'  �#  ,    ='    H3  >�#  d'  7'  �#  ,    T�  �'  ]$  ,   ,   �&   Lk� q�#  U�  |�'  2$   J  W6&  �'  �#  �'   k  J  f%   �'  �#  �'  �#   J�  g7   �'  �#  �'  �#   J?  Ҁ#  (  �#   VpO qO !(  W$   E.  �  $,0  -;  K  :�)  �e  =0  � ?k  "  @�#  �4  AK.  �J  BQ.  �A  O�(  �(  W.   �A  Q�(  �(  W.  ].   �A  V�(  �(  W.  �#   -�
 Y51  _(  �(  �(  c.  w(   -�
 ]�R  k(  )  !)  c.  �(   -� c?  _(  9)  I)  W.  S(  �&   X_ m.   ])  m)  W.  _(  S(   -�3  q89  S(  �)  �)  c.   X.E  ��3  �)  �)  W.  _(  Q.   X�(  ��(  �)  �)  W.  _(   Y_Tp q   G(  ZZD   ��+  [F�   �k   \��   ��"  \�4   �#  \�  � #  (��   �0*  6*  �0   <��   �G*  R*  �0  �0   **   ��}  *  k*  q*  �0   *Ư   �?s  *  �*  �*  �0   *�F   �Ϭ  �0  �*  �*  �0   *�F   ��  �)  �*  �*  �0  �#   *a�   �
�  �0  �*  �*  �0   *a�    ��  �)  +  +  �0  �#   *�:   ,�  *  /+  :+  �0  �)   *�F   		n  �0  S+  ^+  �0  �)   *(*   ��  �)  w+  �+  �0  �)   * I   h�  �0  �+  �+  �0  �)   *�O   7k  �)  �+  �+  �0  �)   *WC   ]�  �0  �+  �+  �0   /{�  k  /�  �   18E  �)  ]*; !1%,  �8  �; N;  �; !v�,  �= !|u.   ^�; !L,  W,  �0  �0   !�  !��= �0  n,  y,  �0  �0   �; !��,  �,  �0   X\ !��: �,  �,  �0   Xf !��8 �,  �,  �0   _�9 !��: �0  �,  �0    %,  (8 !�v-  r< !�%,  �9 !�1   ^(8 !�-  !-  1  1   !�  !�< 1  8-  C-  1  1   )(8 !�S-  ^-  1  1   '8 !�j-  1  �#    �,  �; "/�-  |  "02.   `U  A�.  �-  �1  �#   a��  I�-  �1  �#   `9+  N�.  �-  �1  �#   a��  \�-  �1  �#   b�= !5�-   ,   �� �� W2*  7&.  c8a   dt  d�  �  �  t  d�  dq  d�#  G(  d�)  �)  F  d�  ��  #!�#  �  $ �#  �#  �  ^  �  �  d�  d^  d�  e7   �.  f 3  �  �.  �.  �#  c  d�"  �"  
   du"  u"  /  z"  e�.  /  f e'/  '/  f -/  �.  d"  "  �l  %%   j�  %#%   gtm ,%,�/  ,g  %.�#   �  %/�#  �  %0�#  ��  %1�#  ��  %2�#  ��  %3�#  ��  %4�#  �  %5�#  d�  %6�#   ��  %7%   $~�  %8�#  ( L\�  %>I/  Jѯ  %H6&  	0  >/  >/   J��  %M>/  0  0   T/  J�  %C>/  90  90   >/  J#�  %ak  T0  T0   Z0  T/  J�� %fk  t0  t0   z0  >/  J��  %W0  �0  t0   J[v  %\0  �0  t0   J��  %R,   �0  k  ,   �#  T0   �)  d�0  k  ,  d�)  %,  d�,  d%,  u.  1  d�,  �,  dv-  d�,  h01  i7; "�0   c 1  R�#  B1  j H1  k�5  71  �#  eq  h1  lg%   X1    d #  dz"  d  �.  m�-  �1  nXF  A�1  n\;  A�#  op�T  C�.    m�-  �1  nXF  I�1  n\;  I�#   q�  �1  �1  rh  �1   �.  q�  2  2  rh  �1   m  '2  os__p �]$    q;  52  ?2  rh  ?2   �.  qq  R2  \2  rh  \2   �.  q�  o2  �2  rh  �2  r#  �.   m1  m�-  �2  nXF  N�1  n\;  N�#   q  �2  �2  rh  \2  t__a ��2   o.  q�  �2  �2  rh  �1   qT  �2  3  rh  3  u__n �,  u__c �q   �.  m�  >3  nhR  �>3  nmR  �C3   &.  ,.  q�  V3  `3  rh  \2   q�  n3  �3  rh  \2  t__n �,   q[  �3  �3  rh  �1   m  �3  u__s 9.   m�-  �3  nXF  \�1  n\;  \�#   q  �3  4  rh  4  ov�&  2.  ow__i  0     �.  qy,  4  $4  rh  $4   �0  q�,  74  A4  rh  $4   q�,  O4  Y4  rh  $4   q�  g4  q4  rh  4   x�  q�  �4  �4  rh  4   q�  �4  �4  rh  �4   /  qC-  �4  �4  rh  �4  nF�  !��4   1  1  q^-  �4  �4  rh  �4  r#  �.   y   �5  5  rh  -/   q�  #5  -5  rh  �1   m�  \5  z�e  9.  z�e  9.  u__n 0   q�(  j5  }5  rh  }5  r#  �.   W.  q�  �5  �5  rh  �5  r#  �.   i.  q�(  �5  �5  rh  }5   q}  �5  �5  rh  �5   q�(  �5  �5  rh  }5  �5   ].  q�  6  6  rh  �5  t__a s6   o.  q�  06  :6  rh  �1   y  K6  ^6  rh  ^6  r#  �.   �.  q�  q6  �6  rh  ^6  zv�  k  u__a �6   o.  x#
  q3
  �6  �6  rh  3   q�  �6  �6  rh  3  u__c =q   qy  �6  �6  rh  3  u__s 2�#   q�  7  "7  rh  3  u__s ��#   q�  07  F7  rh  3  u__c �q   q9  T7  g7  rh  3  r#  �.   {a2  ; p$   ��7  �7  |o2  �  {a2  �= �$   ��7  �7  |o2  � }�$&\  ~� �   �   N �7  �7  rh  �7  n�< N�7   �.  �.  {�7  X; �$   �8  s8  |�7  � |�7  ��Y4  �$   P|g4  P��3  �$   ���3  |�3  P��1  �$   d��1  |�1  P    �!  U �8  �8  rh  �7  nm< U�.   {s8  �8 �$   ��8  �8  |�8  � |�8  � q0  �8  �8  rh  3  u__s z�#   qI  �8  9  rh  3  u__s ��#   q�  9  >9  rh  3  u__c -q  ovR'  /E    �o!  z�$�  �X9  �B  �h  �B  ��`�  �B  ��&  |�"  � ��3  �$?   �9  ��3  � ��$?   ��3  � ��$&   ��3  / �%;\     ��6  +%��  �M:  �7  Z �7  ��8  +%��  ���8  Z ��8  ��3  +%   A:  ��3  Z �3%X\   �>%     �"7  >%��  ��;  �97  m �07  �9  >%��  ��#9  m �9  ���  �09  � ��2  >%��  /�:  ��2  ��1  >%   ��2  ��1  >%   -��1     �3  g%   2;  �23  � �'3  "  ��1  k%   3L;  �2  ��1  k%   -��1    �`3  m%��  3�;  �w3  : �n3  X ��&   �w3  z �n3  � �D2  �&   ծ;  �R2   �3  �&	   ׍23  �'3  �    �_%z     ��6  {%��  �Y<  �7  � �7  ��8  {%��  ���8  � ��8  ��3  {%�  M<  ��3  � ��%X\   ��%     � �  �@  s__i �0  �"7  �%8�  ��=  �97  � �07  �9  �%8�  ��#9  � �9  �8�  �09  � ��2  �%   /=  ��2  ��1  �%   ��2  ��1  �%   -��1     �3  �%   29=  �23    �'3  U   ��1  �%   3m=  �2  ��1  �%   -��1    �`3  �%P�  3�=  �w3  m  �n3  �  ��&   �w3  �  �n3  �  �D2  �&   ��=  �R2   �3  �&	   ׍23  �'3  �     ��%z     ��6  �%h�  �z>  �7  �  �7  ��8  �%h�  ���8  �  ��8  ��3  �%��  n>  ��3  �  ��%X\   ��%     �"7  �%��  �@  �97   ! �07  �9  �%��  ��#9   ! �9  ���  �09  "! ��2  �%��  /?  ��2  ��1  �%   ��2  ��1  �%   -��1     �3  &   2E?  �23  @! �'3  h!  ��1  &   3y?  �2  ��1  &   -��1    �`3   &��  3�?  �w3  �! �n3  �! ��&    �w3  �! �n3  �! �D2  �&   ��?  �R2   �3  �&   ׍23  �'3  �!    �&z     ��6  *&��  ��7   " �7  ��8  *&��  ���8   " ��8  ��3  *&�  v@  ��3   " �;&X\   �F&      ��6  p&   ��@  ��6  " ��6  ��8  p&   3��8  " ��8  ��3  p&   }�@  ��3  " �|&X\   ��&    ��6  �&   ~aA  ��6  3" ��6  H" ��2  �&   ?�3  3" ��2  \" ��2  H" ��&�    ��6  �$   |�A  ��6  p" �c6  �$   ���6  �z6  �" �q6  p"   �'6   �B  �T7  ��1  '   #�A  �2  ��1  '   -��1    ��2  
'/   #|�2  ug���2  �" �'   ��2  �" ��2  �" ��2  ' �  ��B  ��2  ��2  # ��1  ' �  V��1  ��1  # � �  ��1  S   �4'.     �$%z   �'p\   �.  m+#  �B  /!T  q  z\C  �	�B  z?)  �	�B   �.  �.  ��!  \@'�  �C  _G  �h  �B  � �?)  \_G  ��8�  JG  ��&  b2.  ## ��B  �'p�  lND  ��B  6# ��B  e# ��2  �'��  �	�C  ��2  e# ��1  �'   ��2  e# ��1  �'   -��1  e#    ��2  �'   �	D  ��2  �# ��1  �'   ��2  �# ��1  �'   -��1  �#    �-5  (   �	�O5  �# �C5  �# �75  �# �(�\    �F7  �'��  l;E  �T7  $ ��1  �'��  #�D  �2  $  ��2  �'��  #��2  4$ ��2  c$ �`(B   ��2  �$ ��2  �$ ��2  `(��  �.E  ��2  �$ ��2  �$ ��1  `(��  V��1  �$ ��1  �$ ���  ��1  %    ��(.     �F7  �'�  l(F  �T7  3% ��1  �'   #yE  �2  3%  ��2  �'(�  #��2  b% ��2  �% �0(0   ��2  �% ��2  �% ��2  0(@�  �F  ��2  �% ��2  & ��1  0(@�  V��1  �% ��1  & �@�  ��1  5&    �J(.     �F7  �(X�  l+G  �T7  U& ��1  �(   #�F  �2  U& ��1  �(   -��1  U&   ��2  �(p�  #��2  w& ��2  �& ��(   ��2  �& ��2  �& ��2  �(��  �G  ��2  ��2  �& ��1  �(��  V��1  ��1  �& ���  ��1  '    ��(.     �z'�\  ��'>9  ��'>9   ��(p\  ��(�\   �.  �2"  ��(�   ��G  �=8 �  � ���  ��&  ��#  ,' �})T#    �q4  =9 �)   ��G  ��)   �{  �)-   ��G  �q4  �)   ֋�)    ��  �)   �q�  H  &H  rh  �4   *  � 6H  zH  rh  4  r#  �.  �ZH  s__i �0   �lH  s__i �0   os__i �0    �&H  �: �)c  ��H  8J  |6H  � ���  BI  �NH  �' �H  *��  �H  �' ��2  *��  �,I  ��2  �' ��2  	( ��1  *��  V��1  �' ��1  	( ���  ��1  (    �+�\  �"+�\    ��  �I  �`H  X( �H  o*(�  �H  �( ��2  o*H�  ��I  ��2  �( ��2  �( ��1  o*H�  V��1  �( ��1  �( �H�  ��1  �(    �+�\  �	+�\  �C+�\    ��*   J  �mH  ��*�\   �A*�\  ��*�\  ��*�\  �8+p\   1!  X HJ  [J  rh  �7  r#  �.   {8J  �= P+6   �vJ  K  |HJ  � �w4  Z+`�  Y��4  �( ��2  Z+��  �J  ��2  ��2  �( ��1  Z+��  V��1  ��1  �( ���  ��1  0)    ���  ��4  C) �y+zH  ��+&\     �L!  q�+W   �3K  RL  �h  �7  � ��< qRL  ��Y4  �+   s�K  �g4  b) ��3  �+   ���3  ��3  b) ��1  �+   d��1  ��1  b)    �w4  �+��  t��4  u) ��2  �+��  'L  ��2  ��2  u) ��1  �+��  V��1  ��1  u) ���  ��1  �)    ��+   ��4  �) ��+zH  ��+&\     �.  �  � gL  �L  rh  4  n< ��L  n4&  �0  ��L  w__i 0   ��L  w__j 0   ��L  w__k 0   ow__l 0  ovR'  O#     2/  {WL  !9 �+�  ��L  �N  |gL  � |pL  �|{L  ����  �M  ��L  �) ��4  c,   ��4  �) ��3  c,   ���3  �) ��3  * ��1  c,   d��1  �) ��1  *     ���  N  ��L  !* ��4  �,   ��4  @* ��3  �,   ���3  S* ��3  g* ��1  �,   d��1  S* ��1  g*     ��,   %N  ��L  |*  � -P   mN  ��L  �
->   ��L  �* �-�\  �)-]  �H--]    �:,]  ��,]  ��,]  �a-�\  �i-zH  �q-K]  �x-�\  ��-p\   �	  7�-�  ��N  �R  �h  4  � ��: 8�.  ���; 8/  ���  �R  v;5 <0  �o8 e�R  �* ��4  �-0�  <�O  �5  �* ��2  �-   ���2  + ��2  + ��1  �-   V��1  + ��1  + ��-   ��1  0+     �H�  �P  �]8 AO#  T+ � : D/  �+ �68 E/  �+ ��9 M/  %, ��; N/  P�`�  &P  �__i G0  h,  � .!   FP  �__l I0  |,  �x�  bP  �__j X0  �,  ��.   �P  �__k Z0  �,  ��-]  �f.]  ��.�\  ��.�\  ��/�\  ��/�\  ��/K]  �0�\   ��4  �.��  d>Q  ��4  �, ��3  �.��  ���3  �, ��3  - ��1  �.��  d��1  �, ��1  -    �H  /��  i�Q  �H  6- ��2  /��  ��Q  ��2  T- ��2  v- ��1  /��  V��1  T- ��1  v- ���  ��1  �-    ��/�\  ��/�\   ���  �__i y0  �- ���  ��; {/  �- �H  S/ �  ~�H  . ��2  S/@�  �{R  ��2  . ��2  Z. ��1  S/@�  V��1  . ��1  Z. �@�  ��1  o.    ��/�\  ��/�\  �0�\      ��/p\  �0p\   �R  d/  ��  , 0`   ��R  �S  �h  4  �. �< -8/  �. ��: -�.  �. �X�  v;5 /0  ��4  10p�  /�S  �5  	/ ��2  70   ���2  3/ ��2  G/ ��1  70   V��1  3/ ��1  G/ �70   ��1  _/     �s0�N  ��0T#    ��  #�0;   ��S  T  �h  4  � �< $8/  ��h8 %'/  �/ ��0�R   m$1  T  op;; $%,    �-  ��0v   �7T  ,U  �h  4  �/ ���  �/  �/ �;5 �0  �/ ���  v�_ ��,  �T  �0��  ��T  ���  �T  �1Q]  �11k]    ��4   1   �U  ��4  0 ��3   1   ���3  *0 ��3  >0 ��1   1   d��1  *0 ��1  >0    ��0~� �   {�4  �(  @1   �GU  �U  |5  � ��2  J1   ���2  S0 ��2  g0 ��1  J1   V��1  S0 ��1  g0 �J1   ��1  0     �D  O�U   _$  ��  P�U  �1  Q�U  ��  W�U   j$  �^  X�U  �U  =V   u$  ��   >V  �B  ?V  ��  E4V   �$  �B   F4V  �C  G4V  �e  H4V  �8  I4V  ��  J4V  �

  X�V   �$  ��  Y�V  ��
  Z�V  ��   `�V  �$  ��  f�V   �$  ��  g�V  ��  h�V  ��  n�V   �$  ��	  o�V  ��  p�V  �H  vW   �$  �`  wW  �w  xW  �   yW  �~  VW   �$  �   �VW  ��  �VW  �  �VW  ��   �VW  ��  �VW  ��	  �VW  ��  ��W   �$  �  ��W  �  ��W  ��  ��W  ��  ��W   �$  ��  ��W  ��  ��W  ��  ��W  �m  �(X   �$  �	  �(X  �2	  �(X  ��  �(X  �9  �(X  �[  �nX   �$  �J  �nX  ��  �nX  �7  �nX  ��  ��X   �$  �I	  ��X  �$	  ��X  ��   ��X   %  �N  ��X  �p  ��X   %  ��  ��X  �:  ��X  ��  ��X  �d   ��X  ��  �8Y   %  �  �8Y  ��  �8Y  ��	  �dY   %%  ��  �dY  �  ؃Y   0%  ��  كY  ��  ڃY  ��  ۃY  �+  �Y   ;%  ��  �Y  ��   �Y  �  ��Y   F%  ��
  ��Y  ��  ��Y  �  �Z   Q%  �   �Z  �F  �Z  ��  �@Z   \%  ��  �@Z  ��  �@Z  ��  3lZ   n%  ��  4lZ  ��   8�Z   y%  ��  9�Z  �l	  =�Z  �%  �N  >�Z  �^  ?�Z  �L  @�Z  �a  D�Z  �%  �B  E�Z  ��	  F�Z  �  G�Z  �  H�Z  �y  I�Z  ��   6[   �%  ��  !6[  ��-   ��  u8 �
	��  9 �
	��  �9 �
	��  �9 �
	��  y= �
	��  B< �
	��  �9 �
	��  �< �
	�[  Gf9 �E�g  H�< �E��  �: �E��  �< �
	�$   ��9 �E�  &�1  ;\  ]$   �mw  ww  �#  X\  �#  �#   �O2  Y2  7   p\  �#   �>  Y  �\  ]$   ���  ��  �#  �\  �&  �&  7    Jww  B�#  �\  �#  �#   �  �\  ]$   ��  ]$  �\  ]$   ��  �e  &�Ӫ  �\  ]$   JY2  Q,   ]  �#   .�  &��  ]$  -]  0   ��d  ]$  K]  ]$  �&  g%   ��  �e= �#  e]  e]   V$  �Y< e]    N   �r   A *B �V  ��       �  (  �  �  �  E   �  �  o  �	  �  qW  !s   int   "�   �  #  .  <h   `  Ds   �  Wh   �  _z   �  es   t   ms   a  us     ~s   �  �s   3  �s   �  �s   H  �s   y  �s     �s   s  �s   T   �s   �  �s   F  �s   �  �s   �  �s     �s   V  �s   3   �  s  N:   �  V:   \	  2s   o  7s   �  <s   �  Cs   �  	s   �  �  3   	
pO qO 
!�  
std  �,  @�  %  0�=  ��  �b  �3   Fe  �s   �#  ��  �&  �q  �3  �=  q  �.  �.   +  eq �<-  �.  �  �.  �.   lt ��1  �.  �  �.  �.   ��  eF  s   �  �.  �.  |   �K  �9  |  �  �.   �(  
!  �.    �.  |  �.   1  �A  �.  6  �.  �.  |   �5  �'  �.  Z  �.  �.  |   �3  �A  �.  ~  �.  |  +   +  :  +  �  �.   6  �C   �P  6  �  �.   �B  $6  �.  �  �.  �.   eof (�:  6  ?  ,N0  6  �.    E  �  9Q  pq  G0  sq   �T  t�  %  {<  B  71   %  �R  ]  71  q   �:  �b;  q  u  {  =1   �T  �4>  �  �  71  �   �T  �QM  �  �  �  =1   �F  ��?  C1  �  �  71  q    I  �O  C1  �  �  71  q   (*  �	H      !  =1  q   �O  �eT    9  D  =1  q   �O  ́?  q  \  g  =1  I1   �$  �   �:  Z�   _� �,   5�.  6�/  7�/  �?  �%   K  \'  �,   �e  _|  �4  c	0  �J  d0  ��  q�  �  '0   ��  s    '0  -0   W  y  '0  s     �  �J  p�  �B  u  �    %  �   !�B  d  D0  �  -0    �e  y�  "[V  �  u   �G  !8   <  x�  �4  {�  �J  |�  �J  N.  `S  �S.  ~J  ��  �J  ��  �%  �%  �K  �u   I  �u  :!  ��/   %H  ��  �   #�3  2�  #�G  7�  #t3  Bn0  $�'  ��O  \0  %V  ��N  �.  ~  �  y0   %3  �o+  �.  �  �  y0   &�P  ��O  �  �  V0   &�M  ��P  �  �  V0   &�,  �-  �  �  V0  u   %�+  ��R  �      V0   %3  �   �  %  5  V0  -0  -0   �/  !�B  V0  Y  u  u  -0   &�O  �|6  l  w  V0  -0   '(  ��6  �  �  V0  -0   (�   �-  �  �  �  V0   )�1  o�*  �  �  V0  -0  u    (�A  $n%  �  �  �  J0   (�A  (�I  �  	  	  P0  �   ("A  ,�%  V0  2	  8	  J0   (�1  2E)  �  P	  V	  J0   (�/  6;&  �  n	  t	  J0   '�>  :�>  �	  �	  P0   (S  A:2  u  �	  �	  J0  u  �   '�#  K�(  �	  �	  J0  u  u  �   (9  S>$  u  �	  
  J0  u  u   (-U  [�7  �.  
  *
  J0  �   *�5  d�-  J
  �  �  u   *	1  m�P  j
  �  �  u   *�3  v\-  �
  �  u  3    *nU  ��-  �
  �  �  �   *nU  �nG  �
  �  �  �   *nU  ��   �
  �  �  �   *nU  �IP  
  �  �  �   �J  �rR  s   )  u  u   '�=  ��H  =  R  P0  u  u  u   'V  �)  f  l  P0   +�'  �D*  \0  ,�0  ��  �  P0   -�0  ��  �  P0  -0   �0  ��  �  P0  b0   �0  ��  �  P0  b0  u  u   �0  ��    P0  b0  u  u  -0   �0  �(  =  P0  �  u  -0   �0  �M  ]  P0  �  -0   �0  �m  �  P0  u  3   -0   ,�0  "�  �  P0  s    .�  *,Q  h0  �  �  P0  b0   .�  2�G  h0  �  �  P0  �   .�  =�%  h0  �  
  P0  3    .S� f�&  �  #  )  P0   .S� q�>  �  B  H  J0   /end y<  �  a  g  P0   /end �6;  �  �  �  J0   .I ��$  �  �  �  P0   .I ��7  �  �  �  J0   .��  �lC  �  �  �  P0   .��  �CM  �  �    J0   .r ��R  u    !  J0   .�K  �r5  u  :  @  J0   .�3  �j=  u  Y  _  J0   0�� �  t  �  P0  u  3    0�� ��F  �  �  P0  u   .I  v  u  �  �  J0   0�E  �|U  �  �  P0  u   0�1  -�  �  �  P0   .�� 5�?  �.      J0   .�:  D�6  �  6  A  J0  u   .�:  UW  �  Z  e  P0  u   /at k
/  �  }  �  J0  u   /at ��7  �  �  �  P0  u   .�F  ��/  h0  �  �  P0  b0   .�F  �k:  h0  �  �  P0  �   .�F  ��H  h0      P0  3    .@  DA:  h0  0  ;  P0  b0   .@  U�1  h0  T  i  P0  b0  u  u   .@  )�D  h0  �  �  P0  �  u   .@  ��*  h0  �  �  P0  �   .@  �6  h0  �  �  P0  u  3    0�G  -aN  �  �  P0  3    �3  �b*  h0    "  P0  b0   .�3  ^ 2  h0  ;  P  P0  b0  u  u   .�3  �=  h0  i  y  P0  �  u   .�3  z�T  h0  �  �  P0  �   .�3  � @  h0  �  �  P0  u  3    0� ��E  �  �  P0  �  u  3    .� �\+  h0  	    P0  u  b0   .� �u>  h0  2  L  P0  u  b0  u  u   .� g|=  h0  e  z  P0  u  �  u   .� "�@  h0  �  �  P0  u  �   .� 9k<  h0  �  �  P0  u  u  3    .� K�'  �  �  �  P0  �  3    .bL  d�R  h0    #  P0  u  u   .bL  t�2  �  <  G  P0  �   .bL  �L&  �  `  p  P0  �  �   .�%  �9F  h0  �  �  P0  u  u  b0   .�%  �|<  h0  �  �  P0  u  u  b0  u  u   .�%  ��T  h0  �  	  P0  u  u  �  u   .�%  ��A  h0  "  7  P0  u  u  �   .�%  b>  h0  P  j  P0  u  u  u  3    .�%  3%  h0  �  �  P0  �  �  b0   .�%  'V7  h0  �  �  P0  �  �  �  u   .�%  <�+  h0  �  �  P0  �  �  �   .�%  Q'S  h0    ,  P0  �  �  u  3    .�%  vj.  h0  E  _  P0  �  �  �  �   .�%  ��9  h0  x  �  P0  �  �  �  �   .�%  �C  h0  �  �  P0  �  �  �  �   .�%  �>/  h0  �  �  P0  �  �  �  �   (�?  ��&  h0    *  P0  u  u  u  3    (�1  �O  h0  B  \  P0  u  u  �  u   ,)  �z-  �  �  u  3   -0   1+E  �3J  �  �  u  3   -0   .�5  ��)  u  �  �  J0  �  u  u   0n	 @D  �  �  P0  h0   .W�  �6  �  
    J0   .�A  %�A  �  )  /  J0   .��  ,Z5  �  H  N  J0   .�(  �;  u  g  |  J0  �  u  u   .�(  I�%  u  �  �  J0  b0  u   .�(  X�5  u  �  �  J0  �  u   .�(  �^   u  �  �  J0  3   u   .�(  v�S  u       J0  b0  u   .�(  	K  u  9  N  J0  �  u  u   .�(  �o?  u  g  w  J0  �  u   .�(  J5  u  �  �  J0  3   u   .NW  ��Q  u  �  �  J0  b0  u   .NW  /�I  u  �  �  J0  �  u  u   .NW  ��,  u       J0  �  u   .NW  ��;  u  9  I  J0  3   u   .�S  ��I  u  b  r  J0  b0  u   .�S  >T?  u  �  �  J0  �  u  u   .�S  05  u  �  �  J0  �  u   .�S  $S:  u  �  �  J0  3   u   .�>  2hL  u      J0  b0  u   .�>  SUB  u  4  I  J0  �  u  u   .�>  Q�2  u  b  r  J0  �  u   .�>  _�K  u  �  �  J0  3   u   .�4  qT  u  �  �  J0  b0  u   .�4  j�K  u  �  �  J0  �  u  u   .�4  ��5  u      J0  �  u   .�4  N.  u  4  D  J0  3   u   .U+  �)  ,  ]  m  J0  u  u   .��  �!1  s   �  �  J0  b0   .��  ��T  s   �  �  J0  u  u  b0   .��  ��O  s   �  �  J0  u  u  b0  u  u   .��  �;.  s       J0  �   .��  ��B  s   4  I  J0  u  u  �   .��  ��,  s   b  |  J0  u  u  �  u   %  !T  3   2�E    2�F  �   3�&  3�7  ,  �o  >8"  �| Cs   4Q  b�   �  4�F c�  4�R  d�  43  e�  4�  f�  4�K  g�  4�@  h�   5all i�  ?6�� ��   :!  ��/    NF  ��0   �E  �|   p0  ��0   �%  ��0  7S  ��0  7�R  ��0  73  ��0  7�$  ��0  7�K  ��0  7�@  ��0  7�@  ��0  '�4  �Z  �  �  0   '�=  y)      0   8��   (  0  �0  |   8�� 8  H  0  �  |   8�� X  c  0  |   8N  s  ~  0  s    8�� �  �  0  �0   '�  �U  �  �  0  �0   (�&  �.  �.  �  �  0   '�F  &�;  �  �  0  �0  �   '�9  )�Q      0  �0  �0   'WR  ,`2  2  B  0  �0  �0   '�S  /=  V  f  0  �0  �0   9e  7,  v  0  �0  |     �$  0   7OD  0  7gP  0  7�F  $�0  3< :id �N    �U  �|   7�I  ��/  '�  �<?  �     �0  �0   ;id �      �0  �0   <id �,   2   �0   =4H  ��(  |  G   �0    �o  u^   d   �0   �o  ~t      �0  �0   -�o  ��   �   �0  �   �o  ��   �   �0  �0  �  �   �o  ��   �   �0  �0  �0  �   5  ��   �   �0  s    �  ��*  �0  !  "!  �0  �0   H�  ��N  ="  :!  @!  �0   U  �9  �.  X!  c!  �0  �0   2  �t*  �.  {!  �!  �0  �0   >jP  �D  �  �!  �0   ?RD  �Q  �0  @�o  7�!  �!  �0  0   A�K  :�N  A�A  =�5  �K  @I  �  �!  �   '�,  CH<  "  ("  �0  �0  �0  �   �  �  1   �  � >,  BW  3�"  C�4  C�$  Cq-  Cc=  Co'  C�5   C�%  � C�8  �CX)  �C�%  �C�  �CaO  �CY=  � CP  �� C�C  ��CwS  �C�O  � C�?  �C�5  �� B
$ g#  C)W  C�   C�U  C�A  C�8  C�P   CEH  �� B�4  �=#  CO   C�7  C(  C�Q  CG  �� B��  �d#  C�R   C�-  C�1  ClO  �� Db4 %  E�N  �=#  E�9  i�"  �P  �H"  F�4  �#  �#  Gdec �#  Ft-  �#  Ghex �#  Fr'  �#  F< �#   Goct �#  @F� �#  �H[)  �#   H�%  "�#   H�  &�#   HdO  )�#   H\=  ,�#   H�P  /�#    H�C  3�#   @FzS  6�#  �F�O  9�#  JH�?  <�#  E�  J#  F�7  N�$  �$  F(  Q�$  F�Q  V�$  FO  Y�$   Gin w�$  z#  Gout z�$   I�M   x%  
,  J�B 1   �b  �3   K:C �1  K�A �1  K�B �1  K�? �1  K�D �1  K_> �1  K]? ��  Fe  �6  �#  �A  �&  �L  LZ  �%  �%  �%  1  s    �= �+D �  �%  �%  1  �0   -H  �C �  &  &  1   V@ �@ 1  &&  6&  1  1  ,   -9  ��<  �%  N&  c&  1  �%  m#  z#   .:H  ?,  �%  |&  �&  1  �%  z#   .X'  F6  s   �&  �&  1   .�D t> ,  �&  �&  1   .!a  *�a  �%  �&  �&  1   .�c  <�c  �%  '  '  1   .�a  R(b  �%  !'  ''  1   .�W  elD ,  @'  P'  1  1  ,   .j> t�B �%  i'  t'  1  "%   .�D �'? �%  �'  �'  1   .�S  �YH  �%  �'  �'  1  "%   .�W  �B  ,  �'  �'  1  %1  ,   "%  ,�B ��'  �'  1   .% ��" 1  (  (  1   .�* �_e  1  4(  :(  1   .�* �e  1  S(  Y(  1   0cb  �Pc  n(  y(  1  s    0��  �R�  �(  �(  1  1  1  1   .� � 1  �(  �(  1   .�-  P  1  �(  �(  1   .�-  �  1  �(   )  1   0� !4  )   )  1  s    0��  +�  5)  E)  1  1  1   M�= @�B %  b)  m)  1  �0   NY@ O�D 1  %  �)  �)  1  1  ,   N09  Z�A �%  %  �)  �)  1  �%  m#  z#   N=H  f> �%  %  �)  *  1  �%  z#   N� s�D s   %  &*  ,*  1   N��  ��? ,  %  M*  S*  1   O�W  -�A ,  %  s*  �*  1  1  ,   N�[  ��C �%  	%  �*  �*  1   Nn\  ��@ �%  
%  �*  �*  1   NZ  �lB �%  %  �*  �*  1  �%   O�W  O`@ ,  %  +  -+  1  %1  ,   NP�  k? �%  %  N+  Y+  1  �%   0�? 2E n+  t+  1   0\b  (a  �+  �+  1  ,   0D tC �+  �+  1  ,   8�B "�+  �+  1  +1   (�  *gE 11  �+  �+  1  +1   �%  !T  3   2�E     %  �>  b�    P�b  3  B,  Q_Tp %   �3  �3   ,  1�;  ��> ,  w,  !T  3   �E    1  1   �U  07  ,  1  1  N    R$   �Y.  �  $,|  -�  K  :I.  �e  =|  � ?�  "  @�  �4  A	0  �J  B0  �A  O-  -  0   �A  Q&-  1-  0  0   �A  VA-  L-  0  s    �
 Y51  �,  d-  o-  !0  �,   �
 ]�R  �,  �-  �-  !0  �,   � c?  �,  �-  �-  0  �,  �   _ m.   �-  �-  0  �,  �,   �3  q89  �,  �-  �-  !0   .E  ��3  .   .  0  �,  0   �(  ��(  4.  ?.  0  �,   Q_Tp 3    �,  3ZD  38E   �� �� �� R2*  7�.  S8   T+  Tq  �  q  +  T�  �  8�/  �{  �   ]�  �  \�   �  �D  !�  �3  "�  U>  #�  &�  $�  �  %�  �*  &�   ڡ  '3   $�U  (3   %TL  )3   &�I  *3   'Q  +3   (�C  ,3   )�J  -3   *1  .�  ,o(  /3   0�U  03   1PL  13   2�I  23   3Q  33   4�C  43   5�J  53   6 P)%  K�  �/  s   �   UGT  P�/  �.  �   s   T3   T�  �,  TI.  I.  �  T'    s   �.  8  �  ,  %  T%  T�  T,  V,   y0  W |  1  �0  �0  �  �  T8"  8"  �  T("  ("  �0  -"  �  V�0  �0  W V�0  �0  W �0  �0  T2"  2"  Xs   1  Y 	1  Z�5  �0  "%  %  
,  �'  T
,  T%    ,  T  T,  [�%  ]1  p1  \h  p1  \#  :0   1  ]W  �1  ^hR  �1  ^mR  �1   �.  �.  ]v  �1  ^hR  ��1  ^mR  ��1   �.  �.  ]~  �1  ___c �1   �.  ]�  �1  ___c  �1   �.  ]�  &2  `hR  $&2  `mR  $+2   �.  �.  a�  [�%  D2  N2  \h  N2   1  [:(  a2  k2  \h  N2   [(  y2  �2  \h  N2   ['  �2  �2  \h  p1  bc�&  T�%    [Y(  �2  �2  \h  p1  ___n �s    [�&  �2  �2  \h  p1  bc�&  >�%    [�'  3  3  \h  N2   [�(  3  #3  \h  N2   [�(  13  ;3  \h  N2   [ )  I3  _3  \h  p1  ___n !s    [B  m3  �3  \h  �3  ^Q  �q   71  T�3  %   ],  �3  Q_Tp %   d__a ¼3  d__b ��3   �3  �3  ]6  �3  `�e  �.  `�e  �.  ___n |   [t+  4  4  \h  p1  ___n ,   [�+  '4  =4  \h  p1  ___n ,   [E)  K4  a4  \h  p1  `ȱ  @a4   �0  e=4  �B `1   ��4  �4  fK4  � fT4  � [m)  �4  �4  \h  p1  1  ,   e�4  �D p1   ��4  �4  f�4  � f�4  �f�4  � [�)  �4  5  \h  p1  �%  m#  z#   e�4  �A �1   �*5  j5  f�4  �f�4  �f5  �f	5  �g_3  �1   \hv3  fm3  �   [�)  x5  �5  \h  p1  �%  z#   ej5  > �1   ��5  �5  fx5  �f�5  �f�5  �g_3  �1   hhv3  fm3  �   [*  �5  �5  \h  p1   e�5  �D �1   �6  6  f�5  �  [,*  )6  36  \h  p1   e6  �? �1   �N6  W6  f)6  �  [�*  e6  o6  \h  p1   eW6  �C �1   ��6  �6  fe6  �  [�*  �6  �6  \h  p1  ___c ��%   e�6  lB �1   ��6  �6  f�6  � f�6  � [-+  �6  7  \h  p1  ___c  �%   e�6  k?  2   �"7  37  f�6  � f�6  � eO1  �? 2   �N7  ]7  i]1  �0 j&2 eO1  DC 02$   �x7  �7  f]1  � kO1  82   Ƣ7  i]1  �0 lG2 mT2�M   n�*  `2�   ��7  �8  oh  p1  � p__s P%1  �0 q__n P,  �rp�  s�&  R,  (1 r��  s�D UB,  h1 k3  �2   U18  i3  �1  t��  �8  s�= XB,  �1 uR'  YB,  v�3  �2��  Z�8  i�3  �1 i�3  �1 i�3  �1 w�2�M   x4  �2   ]y04  i'4  2   r��  z__c b�%  P    [�*  �8  �8  \h  p1  bc�&  ��%  c �  �?0    {�8  �@  3?   �9  �9  f�8  � r �  |�8  %2 }�8  ~k2  .3   �G9  iy2  ]2  ~�1  13   �e9  i�1  |2  g�2  43   ��2  i�2  �2    nS*  @3�   ��9  A;  oh  p1  � p__s .1  �2 q__n .,  �r �  s�&  0,  "3 rH�  s�D 3B,  z3 kk2  `3   3:  iy2  �3  tp�  �:  s�= 6B,  �3 uR'  7B,  v�3  �3��  8g:  i�3  �3 i�3  �3 i�3  4 w�3�M   x�3  �3   ;y4  i4  $4   r��  �__c @�+  74 v�8  w3��  @$;  i�8  U4 r��  |�8  s4 }�8  ~k2  �3   ��:  fy2  S ~�1  4   �;  i�1  �4  g�2  4   ��2  f�2  S   x�1  �3   Ci�1  �4      n�%  4q   �X;  �;  oh  p1  ��ȱ  ��;  �t��  �;  �Y�  Ӭ  � k62  4
   Ӯ;  iD2  �4 l)4 wD4�   ly4 w�4�M   �0  e62  �C �4   ��;  �;  fD2  �l�4 �&  �4#   �<  6<  oh  p1  � q__s �1  �q__n �,  � n6&  �4d   �M<  �<  oh  p1  ��Q  ��%  ��@  �m#  ��^F  �z#  �x�4  5   �i	5  5 i5  /5 i�4  C5 i�4  W5 g_3  5   \iv3  v5 im3  �5    nc&  P5X   ��<  m=  oh  p1  ��j(  �%  ��^F  z#  �gj5  h5   	i�5  �5 y�5  ix5  �5 g_3  h5   hiv3  �5 im3  �5    ��&  �5"   ��=  �=  oh  p1  �  ��&  �54   ��=  �=  oh  p1  � r �  ��&  B,  �5   ��&   6�   ��=  j?  oh  p1  � r �  ��&  ,�%  $6 ��2  (6P�  .?  i�2  i6 �(6   �>  |�2  �6 ~k2  (6   ?[>  iy2  i6  ~S2  +6   ?y>  ia2  �6  g�2  26   Bi�2  7 i�2  *7   rX�  i�2  >7 rX�  }�2  ��8  ]6x�  Ei�8  \7 rx�  |�8  z7 }�8  g�2  �6   ��2  f�2  S      ��2  86��  /i�2  �7 �86   M?  }�2  g�1  <6   Vi�1  �7   r��  i�2  �7 r��  }�2       ��2  �c  �6c   ��?  h@  i�2  8 ��6   �?  |�2  ,8 gk2  �6   ?iy2  ?8   r��  i�2  �8 r��  }�2  ��8  �6��  Ei�8  �8 r��  |�8  �8 }�8  ~�1  �6   �$@  i�1  �8  ~�2  �6   �K@  i�2  9 i�2  )9  gk2  >7   �fy2  S      ��2  (b  P76   ��@  �@  i�2  <9 �T7   �@  |�2  [9 ~k2  T7   U�@  iy2  <9  g�1  \7   Vi�1  n9   r��  i�2  �9 r��  }�2     �''  �7   �A  _A  oh  p1  � �__s e1  ��__n e,  ���7�� � ������  �P'  �7N   �wA  =B  �h  p1  �9 �__c t"%  �9 r�  ��&  v�%  �9 �� w?0  �9 ~k2  �7   w�A  iy2  �:  ~�2  �7   }B  i�2  �: i�2  �:  ~�1  �7   ~ B  i�1  �:  ��1  �70�  zi�1  �:    nt'  �7?   �TB  �B  oh  p1  � rH�  ��&  ��%  ; ~k2  �7   ��B  iy2  ;  ~�2  �7   ��B  i�2  E; i�2  Z;  g�1  8   �i�1  n;    ��'  08B   ��B  �C  �h  p1  �; �__c �"%  �; r`�  ��&  ��%  �; ~3  98   �BC  i3  �;  ~;3  C8   �iC  iR3  �; iI3  �;  ~�1  G8   ��C  i�1  <  ��1  b8��  �f�1  ��_     ��'  �8   ��C  D  oh  p1  � �__s �%1  ��__n �,  ���8�� � ������  [�'  D  &D  \h  p1   eD  �> �8@   �AD  PD  iD  &< j�8 e�2  �" �8   �kD  tD  f3  �  ek2  _e  �8   ��D  �D  fy2  �  eS2  e  �8   ��D  �D  fa2  �  e�2  Pc   9   ��D  �D  f�2  � f�2  � �y(  9   � E  =E  oh  p1  � ��  �1  ��;�  �1  ��P�  �1  � ��(  09   �UE  bE  oh  N2  �  e3  P  @9   �}E  �E  f3  �  e#3  �  P9   ��E  �E  f13  �  e;3  4  `9   ��E  �E  fI3  � fR3  � � )  p9   ��E  F  oh  p1  � �M�  +1  ��u�  +1  � �Y+  �9Z   �3F  �F  �h  p1  G< ~k2  �9   _F  iy2  [<  ~�2  �9   �F  i�2  �< i�2  �<  g�8  �9   i�8  �< ��9   |�8  �< }�8  g�2  �9   �i�2  = i�2  *=     e�3  (a  �9   ��F  	G  f4  � f4  � e4  tC  :   �$G  5G  f'4  � f04  � [�+  CG  YG  \h  p1  `(  "YG   +1  e5G  �@ :E   �yG  �G  iCG  I= iLG  j= jU: ��+  `:   ��G  �G  oh  p1  � ��G  � +1  �G,  p:   �,H  !T  3   �E    ��3  �1  � ��D  �1  ��s:   �Z*  ��.  �ow�:w,    �U  =9H   �   ��   >9H  �B  ?9H  ��  EeH   �   �B   FeH  �C  GeH  �e  HeH  �8  IeH  ��  JeH  �

  X�H   �   ��  Y�H  ��
  Z�H  ��   `�H  �   ��  f�H   �   ��  g�H  ��  h�H  ��  n"I   �   ��	  o"I  ��  p"I  �H  vNI   �   �`  wNI  �w  xNI  �   yNI  �~  �I   �   �   ��I  ��  ��I  �  ��I  ��   ��I  ��  ��I  ��	  ��I  ��  ��I   �   �  ��I  �  ��I  ��  ��I  ��  � J   �   ��  � J  ��  � J  ��  � J  �m  �YJ     �	  �YJ  �2	  �YJ  ��  �YJ  �9  �YJ  �[  ��J     �J  ��J  ��  ��J  �7  ��J  ��  ��J     �I	  ��J  �$	  ��J  ��   �K   "  �N  �K  �p  �#K   -  ��  �#K  �:  �#K  ��  �#K  �d   �#K  ��  �iK   8  �  �iK  ��  �iK  ��	  ѕK   C  ��  ҕK  �  شK   N  ��  ٴK  ��  ڴK  ��  ۴K  �+  ��K   Y  ��  ��K  ��   ��K  �  �L   d  ��
  �L  ��  �L  �  �EL   o  �   �EL  �F  �EL  ��  �qL   z  ��  �qL  ��  �qL  �D  O�L   �  ��  P�L  �1  Q�L  ��  W�L   �  �^  X�L  ��  3�L   �  ��  4�L  ��   8M   �  ��  9M  �l	  =&M  �  �N  >&M  �^  ?&M  �L  @&M  �a  D_M  �  �B  E_M  ��	  F_M  �  G_M  �  H_M  �y  I_M  ��  	 �M   �  ��  	!�M  �  �1  �M  �   ��d  �  �M  �  �  �   �>  Y  N  �   T�.   �L   �{  rG �F �V  ��       (  �  �  �  E   �  �  o  �	  �  qW  !s   int   "�   �  #  .  <h   `  Ds   �  Wh   �  _z   �  es   t   ms   a  us     ~s   �  �s   3  �s   �  �s   H  �s   y  �s     �s   s  �s   T   �s   �  �s   F  �s   �  �s   �  �s     �s   V  �s   3   �  s  	N:   �  	V:   \	  
2s   o  
7s   �  
<s   �  
Cs   �  s   �  �  3   	pO qO !�  
std " �/  @�  ��  Y%+  \%  0a1  vY  �#     _Tp �.  �?  �    �=  �!  �b  �3   Fe  �s   �3  �=  �  �1  �1   e  eq �<-  �1  �  �1  �1   lt ��1  �1  �  �1  �1   ��  eF  s   �  2  2  !   �K  �9  !    2   �(  
!  2  6  2  !  �1   1  �A  2  Z  2  2  !   �5  �'  2  ~  2  2  !   �3  �A  2  �  2  !  e   +  :  e  �  2   p  �C   �P  p  �  �1   �B  $6  �1  �  2  2   eof (�:  p  ?  ,N0  p  2    _� �,   52  6A3  7[3  �?  �%   K  \�  �/   �e  _!  �4  cw3  �J  d}3  ��  q�  �  �3   ��  s�  �  �3  �3   W  y�  �3  s     L  �J  pB  �B    L    %  �   !�B  	  �3  �  �3    �e  y_  "[V  3     �G  !�   <  xL  �4  {k  �J  |w  �J  �1  `S  ��1  ~J  �B  �J  �G  �%  ��  #�K  �   #I  �  #:!  �l3   %H  �~  �   $�3  23  $�G  7�  $t3  B�3  %�'  ��O  �3  &V  ��N  �1  #  )  �3   &3  �o+  �1  @  F  �3   '�P  ��O  Y  _  �3   '�M  ��P  r  x  �3   '�,  �-  �  �  �3     &�+  ��R  �  �  �  �3   &3  �   �  �  �  �3  �3  �3   �/  !�B  �3  �      �3   '�O  �|6      �3  �3   ((  ��6  0  ;  �3  �3   )�   �-  �  S  Y  �3   *�1  o�*  �  m  �3  �3      )�A  $n%  �  �  �  �3   )�A  (�I  �  �  �  �3  �   )"A  ,�%  �3  �  �  �3   )�1  2E)  i  �  �  �3   )�/  6;&  i      �3   (�>  :�>  -  3  �3   )S  A:2    K  [  �3    �   (�#  K�(  o  �  �3      �   )9  S>$    �  �  �3       )-U  [�7  �1  �  �  �3  �   +�5  d�-  �  �  �     +	1  m�P  	  �  �     +�3  v\-  /	  �    3    +nU  ��-  O	  �  i  i   +nU  �nG  o	  �  u  u   +nU  ��   �	  �  �  �   +nU  �IP  �	  �  �  �   �J  �rR  s   �	       (�=  ��H  �	  �	  �3         (V  �)  
  
  �3   ,�'  �D*  �3  -�0  �2
  8
  �3   .�0  �H
  S
  �3  �3   �0  �c
  n
  �3  �3   �0  �~
  �
  �3  �3       �0  ��
  �
  �3  �3      �3   �0  ��
  �
  �3  �    �3   �0  ��
    �3  �  �3   �0  �  '  �3    3   �3   -�0  "8  C  �3  s    /�  *,Q  �3  \  g  �3  �3   /�  2�G  �3  �  �  �3  �   /�  =�%  �3  �  �  �3  3    /S� f�&  i  �  �  �3   /S� q�>  u  �  �  �3   0end y<  i      �3   0end �6;  u  %  +  �3   /I ��$  �  D  J  �3   /I ��7  �  c  i  �3   /��  �lC  �  �  �  �3   /��  �CM  �  �  �  �3   /r ��R    �  �  �3   /�K  �r5    �  �  �3   /�3  �j=    �    �3   1�� �    )  �3    3    1�� ��F  >  I  �3     /I  v    b  h  �3   1�E  �|U  }  �  �3     1�1  -�  �  �  �3   /�� 5�?  �1  �  �  �3   /�:  D�6  ]  �  �  �3     /�:  UW  Q  �  
  �3     0at k
/  ]  "  -  �3     0at ��7  Q  E  P  �3     /�F  ��/  �3  i  t  �3  �3   /�F  �k:  �3  �  �  �3  �   /�F  ��H  �3  �  �  �3  3    /@  DA:  �3  �  �  �3  �3   /@  U�1  �3  �    �3  �3       /@  )�D  �3  '  7  �3  �     /@  ��*  �3  P  [  �3  �   /@  �6  �3  t  �  �3    3    1�G  -aN  �  �  �3  3    2�3  �b*  �3  �  �  �3  �3   /�3  ^ 2  �3  �  �  �3  �3       /�3  �=  �3      �3  �     /�3  z�T  �3  7  B  �3  �   /�3  � @  �3  [  k  �3    3    1� ��E  �  �  �3  i    3    /� �\+  �3  �  �  �3    �3   /� �u>  �3  �  �  �3    �3       /� g|=  �3  
    �3    �     /� "�@  �3  8  H  �3    �   /� 9k<  �3  a  v  �3      3    /� K�'  i  �  �  �3  i  3    /bL  d�R  �3  �  �  �3       /bL  t�2  i  �  �  �3  i   /bL  �L&  i      �3  i  i   /�%  �9F  �3  .  C  �3      �3   /�%  �|<  �3  \  {  �3      �3       /�%  ��T  �3  �  �  �3      �     /�%  ��A  �3  �  �  �3      �   /�%  b>  �3  �    �3        3    /�%  3%  �3  (  =  �3  i  i  �3   /�%  'V7  �3  V  p  �3  i  i  �     /�%  <�+  �3  �  �  �3  i  i  �   /�%  Q'S  �3  �  �  �3  i  i    3    /�%  vj.  �3  �    �3  i  i  �  �   /�%  ��9  �3    7  �3  i  i  �  �   /�%  �C  �3  P  j  �3  i  i  i  i   /�%  �>/  �3  �  �  �3  i  i  u  u   )�?  ��&  �3  �  �  �3        3    )�1  �O  �3  �    �3      �     ,)  �z-  �  %    3   �3   3+E  �3J  �  H    3   �3   /�5  ��)    a  v  �3  �       1n	 @D  �  �  �3  �3   /W�  �6  �  �  �  �3   /�A  %�A  �  �  �  �3   /��  ,Z5  E  �  �  �3   /�(  �;      !  �3  �       /�(  I�%    :  J  �3  �3     /�(  X�5    c  s  �3  �     /�(  �^     �  �  �3  3      /�(  v�S    �  �  �3  �3     /�(  	K    �  �  �3  �       /�(  �o?        �3  �     /�(  J5    5  E  �3  3      /NW  ��Q    ^  n  �3  �3     /NW  /�I    �  �  �3  �       /NW  ��,    �  �  �3  �     /NW  ��;    �  �  �3  3      /�S  ��I        �3  �3     /�S  >T?    0  E  �3  �       /�S  05    ^  n  �3  �     /�S  $S:    �  �  �3  3      /�>  2hL    �  �  �3  �3     /�>  SUB    �  �  �3  �       /�>  Q�2        �3  �     /�>  _�K    0  @  �3  3      /�4  qT    Y  i  �3  �3     /�4  j�K    �  �  �3  �       /�4  ��5    �  �  �3  �     /�4  N.    �  �  �3  3      /U+  �)  �      �3       /��  �!1  s   +  6  �3  �3   /��  ��T  s   O  d  �3      �3   /��  ��O  s   }  �  �3      �3       /��  �;.  s   �  �  �3  �   /��  ��B  s   �  �  �3      �   /��  ��,  s     !  �3      �     �  !T  3   4�E  Y  4�F  L   5�&  5�7  �  �o  >�   �| Cs   6Q  bv   ]  6�F cv  6�R  dv  63  ev  6�  fv  6�K  gv  6�@  hv   7all iv  ?8�� �,   :!  �l3    NF  �"4   �E  �!   p0  �"4   �%  �.4  9S  �44  9�R  �44  93  �44  9�$  �44  9�K  �44  9�@  �44  9�@  �?4  (�4  �Z  �  �  �3   (�=  y)  �  �  �3   :�� �  �  �3  U4  !   :�� �  �  �3  �  !   :�� �    �3  !   :N    #  �3  s    :�� 3  >  �3  U4   (�  �U  R  ]  �3  U4   )�&  �.  �1  u  {  �3   (�F  &�;  �  �  �3  [4  ]   (�9  )�Q  �  �  �3  [4  J4   (WR  ,`2  �  �  �3  [4  4   (�S  /=  �    �3  4  (4   ;e  7,    �3  (4  !     �$  �3   9OD  �3  9gP  �3  9�F  $�3  5< <id ��   �U  �!   9�I  �l3  (�  �<?  �  �  4  4   =id ��  �  4  4   >id ��  �  4   ?4H  ��(  !  �  4    �o  u  	  �3   �o  ~  $  �3  4   .�o  �4  ?  �3  �   �o  �O  d  �3  4  �  ]   �o  �t  �  �3  4  4  ]   5  ��  �  �3  s    2�  ��*  4  �  �  �3  4   2H�  ��N  �   �  �  
4   2U  �9  �1  �     
4  4   22  �t*  �1      +   
4  4   @jP  �D  Q  F   4   ARD  �Q  4  B�o  7g   r   �3  �3   C�K  :�N  C�A  =�5  �K  @I  ]  �   ]   (�,  CH<  �   �   �3  4  4  ]   b  ]  �   Q  � >�  DW  3|!  E�4  E�$  Eq-  Ec=  Eo'  E�5   E�%  � E�8  �EX)  �E�%  �E�  �EaO  �EY=  � EP  �� E�C  ��EwS  �E�O  � E�?  �E�5  �� D
$ g�!  E)W  E�   E�U  E�A  E�8  E�P   EEH  �� D�4  ��!  EO   E�7  E(  E�Q  EG  �� Fb4 �%  G�3 �"  E�3  Ex0 EC5  H�3 ��"   '5 �a4    � ��"   �U  �s    :!  �l3  :�3 �^"  s"  a4  �"  s   a4   (�4  ��2 �"  �"  a4   *�=  �]- s   �"  a4    I>. �g4  H�4 ��"   ?6 ��    �+ �%   !�4 ��"  �4    J�#  E�0  I�  J�!  /n4 '�T  -#  '#  -#  �5   �P  ��   /n4 2�t  -#  R#  ]#  �5  -#   /�/ m��  �,  v#  |#  �5   /�/ v2  �,  �#  �#  �5  �,   /l6 ��K  �,  �#  �#  �5   /l6 �6N  �,  �#  �#  �5  �,   /-H  ��`  Q  �#  $  �5   K�4  $  -#  Ldec $  Kt-  $  Lhex $  Kr'  $  K< $   Loct $  @K� $  �M[)  $   M�%  "$   M�  &$   MdO  )$   M\=  ,$   M�P  /$    M�C  3$   @KzS  6$  �K�O  9$  JM�?  <$  K�7  N%  #  K(  Q%  K�Q  V%  KO  Y%   I�9  i|!  Lin wb%  H%  Lout zb%  /�= ��, Q  �%  �%  �5  4   Nf3 �, �%  �5    �!  O�E  �B�!  �)  �!   P I _�4  p�b  K3   PXF `�%  tP�F a�1  uPH b�4  xb  V5*  P�F e�4  |&  '<  X+  PH g�4  �+&  F Z(+  PjF i�4  �I&  2}F sQI �  &  �&  �4   2`F w'I �1  �&  �&  �4   2�M  ��B  #  �&  �&  �4   Q�1  )�%  �&  �&  �4  #   QeU  ��4  �&  �&  �4  #   QbU  �IQ  '  '  �4  #   2�=  �93  �1  6'  <'  �4   Reof �RH �1  T'  Z'  �4   2Z  �4O  �1  r'  x'  �4   Rbad �&H �1  �'  �'  �4   29U  ؍0  #  �'  �'  �4   Q9U  ��H �'  �'  �4  #   SaV  �'  �'  �4  �4   T`V  �%  (  (  �4  s    0tie !�G  �4  )(  /(  �4   0tie -��  �4  H(  S(  �4  �4   /3F  ;�S  �4  l(  r(  �4   23F  5u�  �4  �(  �(  �4  �4   2uF ?�E �4  �(  �(  �4  �4   /[F l�L  �%  �(  �(  �4   /[F ��@  �%  �(  �(  �4  �%   2�= r�H Q  )  )  �4  4   /g�  �(F 3   7)  G)  �4  �%  3    /��  ��$  �%  `)  k)  �4  3    -aV  �|)  �)  �4   Qi3 ~P4  �)  �)  �4  �4   Q�G ��E �)  �)  �4  4   !T  3   4�E  Y   5�8  F�M  5*  2-H  �C Q  �)  �)  S5   2�= �+D Q  *  "*  �4  4   !T  3   4�E  Y   F�+  +  /��  a�)  b*  W*  b*  �6  3    I�b  �3   /g�  ��  3   �*  �*  �6  b*  3    UKC  3�T  b*  5*  �*  �*  �6  3    U҉  d�  3   5*  �*  �*  �6  b*  3    ;+3  ��3  +  �6    F"(  (+  !T  3   4QJ  I+   F�p  D+  !T  3   4�  �,   �%  ;G  آ,  /   }'  ��)  #(T  ��4   #�U  ��1  �E  ��)  "  ��+  �+  �4  �4   "  ��+  �+  �4  �4   2�  �'V  �4  �+  �+  �4  3    /*  )A  �4  �+  ,  �4   /�F  	j8  �4  ,  (,  �4  s    /�F  �8  �4  A,  G,  �4   /V  �0  �1  `,  f,  �4   /�E  L  �4  ,  �,  �4  �  �,   !T  3   �E  Y   I+  �>  bA  ��  v�,  �#    V_Tp 3   �.  �   �?  �  �   w3   ��  2b.  �,   }'  C�)  #(T  a�4   Fe  Bp  #�>  b-  �b  @3   (� Db.  X�  fW-  ]-  �4   X�  pm-  x-  �4  �4   X�  t�-  �-  �4  �4   2*  {p  /-  �-  �-  �4   2�F  �C�  �4  �-  �-  �4   2�F  �ޙ  �,  �-  �-  �4  s    2|�  ���  �1  
.  .  �4   5   &  �%�  -  ,.  2.  �4   &��  Ú�  �1  I.  O.  �4   !T  3   �E  Y   5�Y  �,  �)  W�*  ��!  �.  �!  �!   5*  W*  ��!  �.  �!  �!   W	W  �17  �.  77  �!   �!  WN  .�7  �.  �R  5*  �6   t4 _�/ �.  �   X	@  8�N  3/�  h��  �1  )/  �R  5*  4   3}`  ��d  �7  K/  �R  5*  4   3�g  hL�  �1  m/  �R  +  4   3��  �Ҁ  �L  �/  �R  +  4   +  39�  h|�  �1  �/  �R  (+  4   3c�  ��w  �L  �/  �R  (+  4   (+   Y$   ��1  �  $,!  -A  K  :�1  �e  =!  � ?�  "  @�  �4  Aw3  �J  B}3  �A  OV0  \0  �3   �A  Ql0  w0  �3  �3   �A  V�0  �0  �3  s    2�
 Y51  0  �0  �0  �3  .0   2�
 ]�R  "0  �0  �0  �3  :0   2� c?  0  �0   1  �3  
0  �   Q_ m.   1  $1  �3  0  
0   2�3  q89  
0  <1  B1  �3   Q.E  ��3  V1  f1  �3  0  }3   Q�(  ��(  z1  �1  �3  0   V_Tp 3    �/  5ZD  58E  Z��  I�1  5  s    [��  \5  s     �� �� �� Y2*  7�1  \8(   ]e  ]�  �  �  e  ]�  �  8A3  #�{  �   #]�  �  #\�   �  #�D  !�  #�3  "�  #U>  #�  #&�  $�  #�  %�  #�*  &�   #ڡ  '3   $#�U  (3   %#TL  )3   &#�I  *3   '#Q  +3   (#�C  ,3   )#�J  -3   *#1  .�  ,#o(  /3   0#�U  03   1#PL  13   2#�I  23   3#Q  33   4#�C  43   5#�J  53   6 W)%  K�  [3  s   �   ^GT  Pf3  2  �    s   ]3   ]�  �/  ]�1  �1  L  ]�    s   �  L  �  �  ]�  ]L  ]�  _,   �3  ` !  �  �3  �3  �  Q  ]�   �   b  ]�   �   (4  �   �  _4  ?4  ` _J4  J4  ` P4  4  ]�   �   "  m4  a�4  �!  �4  s    ]�!  �"  �)  �)  &&  D&  b&  D+  �%  ]�%  ]D+  \+  I+  ]�+  ]I+  �,  �,  �,  ];-  g.  ]�,  ]g.  l3  b�1  -5  cXF  I5  c\;  Is    d�'  ;5  N5  eh  N5  e#  �3   �4  l.  d�)  g5  q5  eh  q5   S5  bq.  �5  f__a ��!  f__b ��!   b�1  �5  cXF  \5  c\;  \s    �%  d#  �5  �5  eh  �5   �5  �!  d9#  �5  6  eh  6  g�%  2-#  hi'U  4-#    �5  d]#  &6  06  eh  �5   d|#  >6  b6  eh  6  g�6  v�,  hi'U  x�,    d�#  p6  z6  eh  �5   d�#  �6  �6  eh  6  g�R  ��,  hi'U  ��,    �.  d>*  �6  �6  eh  �6  j__c a3    �6  d�&  �6  �6  eh  �6   �4  b�.  7  f__a ��!  f__b ��!   dZ'  '7  17  eh  �6   ]�.  ]�!  b�.  ^7  f__a �^7  f__b ��!   77  d�'  q7  {7  eh  �6   dS(  �7  �7  eh  �6   d�#  �7  �7  eh  �5   ]�.  b�.  �7  �R  5*  f__f .�6   do*  �7  8  eh  �6  j__c �b*  g�  �3   hk__t ��    d�(  8  &8  eh  �6   d�"  48  >8  eh  >8   �4  ds"  Q8  [8  eh  [8   a4  d(  n8  x8  eh  �6   d/(  �8  �8  eh  N5  gl�  -�4  hi'U  /�4    d�'  �8  �8  eh  N5  cF �#   d�*  �8  �8  eh  �6  j__c 33    l�8  �T  ��   �9  9  m�8  � m�8  � d�*  +9  M9  eh  �6  j__c db*  g�  d3    l9  �  ��   �h9  �9  m+9  � m49  �m@9  � l-5  ~H �:   ��9  �9  m;5  � n�:o� �   l-5  �F �:!   ��9  :  m;5  � p-5  �:   �9  q;5  �= r�: s�:�L   tg&  �:   �:  ':  uh  �6  �  t�&  �:   �>:  c:  uh  �6  � v7  �:   xm'7  �   l�6  �B   ;   �~:  �:  m�6  �  t�&  ;2   ��:  �:  uh  N5  � w�%  )#  �xv5  0;   .�:  q�5  �= q�5  �=  yB;�.   t�&  P;   ��:  S;  uh  N5  � z�%  �#  �= xv5  T;   �@;  q�5  �= q�5  >  {d;�:  o� �   t�&  p;   �j;  �;  uh  N5  � w�%  �#  �x=7  {;   ��;  qR7  > qG7  ;> vv5  {;   �q�5  > q�5  `>   y�;�L   t'  �;   ��;  �;  uh  �6  �  t<'  �;   �<  <  uh  �6  �  l7  4O  �;   �9<  B<  m'7  �  tx'  �;   �Y<  f<  uh  �6  �  lc7  �0  �;   ��<  �<  mq7  �  l�8  �H �;   ��<  �<  m�8  � q�8  t> {�;�:  o� �   l`8  �G   <   ��<  �<  mn8  �  lx8  ��  <   �=  *=  m�8  � m�8  �|<
   }�8  P  l{7  �S   <   �E=  N=  m�7  �  tr(  0<!   �e=  �=  uh  N5  � w(  5�4  �|8<   ~'U  7�4  �> yJ<�:    dG)  �=  �=  eh  �6  j__c �3    8  �L  `<p   ��=  }>  m8  � ��=  �<�  p��=   q�=  �> ��7  �<(�  �2>  q�7  �> y�<�.   ��6  �<@�  �q�6  �> q�6  ? |�<+   q�6  !? q�6  6? y�<�*      d�(  �>  �>  eh  N5  g�R  ��%  hi'U  ��%    }>  �@  �<|   ��>  �?  m�>  � m�>  ��X�  ��>  I? �8  �<x�  �q8  g? ��=  �<��  p��=   q�=  �? ��7  �<��  �M?  q�7  �? yL=�.   ��6  �<��  �q�6  �? q�6  @ |=3   q�6  #@ q�6  8@ y=�*        �)  P=�   ��?  E@  uh  �6  � �__c ��%  ���  �3   ���7  e=��  �@  q�7  K@ y�=�.   ��7  i=��  �q�7  t@ q�7  �@ q�7  "A ���  � 8  KA    ��=  �$  �=b   �a@  �@  m�=  � m�=  ���7  �=�  ��@  q�7  iA yB>�.   ��6  �=0�  �q�6  �A q�6  �A �P�  q�6  B q�6  &B y>�*     dk)  �@  �@  eh  N5   l�@  �F P>J   �A  !A  m�@  � r^> t�)  �>�   �8A  �A  uh  N5  � wȱ  ��A  �y�>/  y�>)/  y�>K/  y�>m/  y�>�/  y?�/  y0?K/  yS?�/   4  d�)  �A  �A  eh  �A  cȱ  ��A  h�Y�  �Q    �4  4  ��(  p?�   ��A  �B  uh  N5  �wȱ  r�B  ��h�  �B  �'U  tQ  � x�7  �?   tIB  q�7  EB r�? x{7  �?   wfB  q�7  qB  ��A  �?��  x�B  q�A  �B q�A  �B ���  ��A  xY5  �?   ӺB  qg5  �B r�? y�?�  r�?  y�?u%  r�?y�?!A  r�?r@ y@�L   4  t�)   @H   �C  ?C  uh  N5  � w(  ~�4  �y3@�%  y?@!A   d�'  MC  cC  eh  N5  g(  �4   l?C  0G p@p   �~C  �C  mMC  � mVC  �r�@y�@�B  r�@y�@�L   ��(  �@_  ��C  �F  uh  N5  Sw?)  ?�F  U���  �3 I�4  V��1 Ma4  WxC8  A   OQD  �Q8  ��5  A   ���5  ��5  v5  A   d�!5  �5     ���  jD  �__i Zs   R �8  �A��  c�D  �8  ��=  �B��  p��=  ��=  ��7  �B�  ��D  ��7   ��6  �B0�  ���6  ��6  |�B4   ��6  ��6      x�5  �A   _#E  ��5  ��5  |�A   �6    xz6  �A   `SE  ��6  ��6  |�A   ��6    x06  �A   a�E  �>6  �G6  |�A   �T6    x`8  �A   b�E  �n8   xx8  �A   b�E  ��8  ��8  |�A   ��8    �}>  �AH�  c�F  ��>  ��>  �H�  ��>  �8  �Ap�  ��8  ��=  �B��  p��=  ��=  p�7  �B   �HF  ��7   ��6  �B��  ���6  ��6  |C6   ��6  ��6        ��7  �A��  d�F  ��7   xc7  �A   j�F  �q7   x�8  �A   j�F  ��8  ��8   v&8  PB   I�48     �4  �U  =�F   �   ��   >�F  �B  ?�F  ��  E+G   �   �B   F+G  �C  G+G  �e  H+G  �8  I+G  ��  J+G  �

  X~G   �   ��  Y~G  ��
  Z~G  ��   `�G  �   ��  f�G   �   ��  g�G  ��  h�G  ��  n�G   �   ��	  o�G  ��  p�G  �H  vH   �   �`  wH  �w  xH  �   yH  �~  MH   �   �   �MH  ��  �MH  �  �MH  ��   �MH  ��  �MH  ��	  �MH  ��  ��H   �   �  ��H  �  ��H  ��  ��H  ��  ��H   �   ��  ��H  ��  ��H  ��  ��H  �m  �I     �	  �I  �2	  �I  ��  �I  �9  �I  �[  �eI     �J  �eI  ��  �eI  �7  �eI  ��  ��I     �I	  ��I  �$	  ��I  ��   ��I   "  �N  ��I  �p  ��I   -  ��  ��I  �:  ��I  ��  ��I  �d   ��I  ��  �/J   8  �  �/J  ��  �/J  ��	  �[J   C  ��  �[J  �  �zJ   N  ��  �zJ  ��  �zJ  ��  �zJ  �+  �J   Y  ��  �J  ��   �J  �  ��J   d  ��
  ��J  ��  ��J  �  �K   o  �   �K  �F  �K  ��  �7K   z  ��  �7K  ��  �7K  �D  	OcK   �  ��  	PcK  �1  	QcK  ��  	W�K   �  �^  	X�K  ��  
3�K   �  ��  
4�K  ��   
8�K   �  ��  
9�K  �l	  
=�K  �  �N  
>�K  �^  
?�K  �L  
@�K  �a  
D%L  �  �B  
E%L  ��	  
F%L  �  
G%L  �  
H%L  �y  
I%L  ��   xL   �  ��  !xL  �  !�1  �L  �   ��  ]�/  ]�/  �>  Y  �    [8   ��  MJ M �V  @�      � (  _� �7   �  �  8k  �{  k   ]�  k  \�   k  �D  !k  �3  "k  U>  #k  &�  $k  �  %k  �*  &k   ڡ  'q  $�U  (q  %TL  )q  &�I  *q  'Q  +q  (�C  ,q  )�J  -q  *1  .k  ,o(  /q  0�U  0q  1PL  1q  2�I  2q  3Q  3q  4�C  4q  5�J  5q  6 q  �  std   -$  5>   6-$  7Y$  @&  	%  0�=  �n  �b  �q  Fe  �G$  
�3  �=  �  &*  ,*   �  eq �<-  2*    ,*  ,*   lt ��1  2*  !  ,*  ,*   ��  eF  G$  E  9*  9*  n   �K  �9  n  _  9*   �(  
!  9*  �  9*  n  ,*   1  �A  ?*  �  ?*  9*  n   �5  �'  ?*  �  ?*  9*  n   �3  �A  ?*  �  ?*  n  �   +  :  �  	  E*   �  �C   �P  �  (  ,*   �B  $6  2*  G  E*  E*   eof (�:  �  ?  ,N0  �  E*    _� 	�7   �?  	�%   K  
\  >&   �e  
_n  �4  
cK*  �J  
dQ*  ��  
q�  �  i*   ��  
s�  �  i*  o*   W  
y�  i*  G$    �  �J  pz  �B  R  �   %  k   �B  A  �*  k  o*    �e  y�  [V  k  R  �G  !   <  x�  �4  {�  �J  |�  �J  �'  `S  ��)  ~J  �z  �J  �  �%  �  �K  �R   I  �R  :!  �|*   %H  ��  �   �3  2k  �G  7T$  t3  B�*  �'  ��O  �*  V  ��N  2*  [  a  �*   3  �o+  2*  x  ~  �*   �P  ��O  �  �  �*   �M  ��P  �  �  �*   �,  �-  �  �  �*  R   �+  ��R  k  �  �  �*   3  �   k      �*  o*  o*   �/  !�B  �*  6  R  R  o*   �O  �|6  I  T  �*  o*    (  ��6  h  s  �*  o*   !�   �-  k  �  �  �*   "�1  o�*  k  �  �*  o*  R    !�A  $n%  k  �  �  �*   !�A  (�I  k  �  �  �*  k   !"A  ,�%  �*      �*   !�1  2E)  �  -  3  �*   !�/  6;&  �  K  Q  �*    �>  :�>  e  k  �*   !S  A:2  R  �  �  �*  R  N$    �#  K�(  �  �  �*  R  R  N$   !9  S>$  R  �  �  �*  R  R   !-U  [�7  2*  �    �*  N$   #�5  d�-  '  k  N$  R   #	1  m�P  G  k  N$  R   #�3  v\-  g  k  R  q   #nU  ��-  �  k  �  �   #nU  �nG  �  k  �  �   #nU  ��   �  k  k  k   #nU  �IP  �  k  N$  N$   �J  �rR  G$  	  R  R    �=  ��H  	  /	  �*  R  R  R    V  �)  C	  I	  �*   $�'  �D*  �*  %�0  �j	  p	  �*   &�0  ��	  �	  �*  o*   �0  ��	  �	  �*  �*   �0  ��	  �	  �*  �*  R  R   �0  ��	  �	  �*  �*  R  R  o*   �0  �
  
  �*  N$  R  o*   �0  �*
  :
  �*  N$  o*   �0  �J
  _
  �*  R  q  o*   %�0  "p
  {
  �*  G$   '�  *,Q  �*  �
  �
  �*  �*   '�  2�G  �*  �
  �
  �*  N$   '�  =�%  �*  �
  �
  �*  q   'S� f�&  �       �*   'S� q�>  �    %  �*   (end y<  �  >  D  �*   (end �6;  �  ]  c  �*   'I ��$  �  |  �  �*   'I ��7  �  �  �  �*   '��  �lC  �  �  �  �*   '��  �CM  �  �  �  �*   'r ��R  R  �  �  �*   '�K  �r5  R      �*   '�3  �j=  R  6  <  �*   )�� �  Q  a  �*  R  q   )�� ��F  v  �  �*  R   'I  v  R  �  �  �*   )�E  �|U  �  �  �*  R   )�1  -�  �  �  �*   '�� 5�?  2*  �  �  �*   '�:  D�6  �      �*  R   '�:  UW  �  7  B  �*  R   (at k
/  �  Z  e  �*  R   (at ��7  �  }  �  �*  R   '�F  ��/  �*  �  �  �*  �*   '�F  �k:  �*  �  �  �*  N$   '�F  ��H  �*  �  �  �*  q   '@  DA:  �*      �*  �*   '@  U�1  �*  1  F  �*  �*  R  R   '@  )�D  �*  _  o  �*  N$  R   '@  ��*  �*  �  �  �*  N$   '@  �6  �*  �  �  �*  R  q   )�G  -aN  �  �  �*  q   *�3  �b*  �*  �  �  �*  �*   '�3  ^ 2  �*    -  �*  �*  R  R   '�3  �=  �*  F  V  �*  N$  R   '�3  z�T  �*  o  z  �*  N$   '�3  � @  �*  �  �  �*  R  q   )� ��E  �  �  �*  �  R  q   '� �\+  �*  �  �  �*  R  �*   '� �u>  �*    )  �*  R  �*  R  R   '� g|=  �*  B  W  �*  R  N$  R   '� "�@  �*  p  �  �*  R  N$   '� 9k<  �*  �  �  �*  R  R  q   '� K�'  �  �  �  �*  �  q   'bL  d�R  �*  �     �*  R  R   'bL  t�2  �    $  �*  �   'bL  �L&  �  =  M  �*  �  �   '�%  �9F  �*  f  {  �*  R  R  �*   '�%  �|<  �*  �  �  �*  R  R  �*  R  R   '�%  ��T  �*  �  �  �*  R  R  N$  R   '�%  ��A  �*  �    �*  R  R  N$   '�%  b>  �*  -  G  �*  R  R  R  q   '�%  3%  �*  `  u  �*  �  �  �*   '�%  'V7  �*  �  �  �*  �  �  N$  R   '�%  <�+  �*  �  �  �*  �  �  N$   '�%  Q'S  �*  �  	  �*  �  �  R  q   '�%  vj.  �*  "  <  �*  �  �  k  k   '�%  ��9  �*  U  o  �*  �  �  N$  N$   '�%  �C  �*  �  �  �*  �  �  �  �   '�%  �>/  �*  �  �  �*  �  �  �  �   !�?  ��&  �*  �    �*  R  R  R  q   !�1  �O  �*    9  �*  R  R  N$  R   ,)  �z-  k  ]  R  q  o*   ++E  �3J  k  �  R  q  o*   '�5  ��)  R  �  �  �*  k  R  R   )n	 @D  �  �  �*  �*   'W�  �6  N$  �  �  �*   '�A  %�A  N$      �*   '��  ,Z5  }  %  +  �*   '�(  �;  R  D  Y  �*  N$  R  R   '�(  I�%  R  r  �  �*  �*  R   '�(  X�5  R  �  �  �*  N$  R   '�(  �^   R  �  �  �*  q  R   '�(  v�S  R  �  �  �*  �*  R   '�(  	K  R    +  �*  N$  R  R   '�(  �o?  R  D  T  �*  N$  R   '�(  J5  R  m  }  �*  q  R   'NW  ��Q  R  �  �  �*  �*  R   'NW  /�I  R  �  �  �*  N$  R  R   'NW  ��,  R  �  �  �*  N$  R   'NW  ��;  R    &  �*  q  R   '�S  ��I  R  ?  O  �*  �*  R   '�S  >T?  R  h  }  �*  N$  R  R   '�S  05  R  �  �  �*  N$  R   '�S  $S:  R  �  �  �*  q  R   '�>  2hL  R  �  �  �*  �*  R   '�>  SUB  R    &  �*  N$  R  R   '�>  Q�2  R  ?  O  �*  N$  R   '�>  _�K  R  h  x  �*  q  R   '�4  qT  R  �  �  �*  �*  R   '�4  j�K  R  �  �  �*  N$  R  R   '�4  ��5  R  �  �  �*  N$  R   '�4  N.  R    !  �*  q  R   'U+  �)  	  :  J  �*  R  R   '��  �!1  G$  c  n  �*  �*   '��  ��T  G$  �  �  �*  R  R  �*   '��  ��O  G$  �  �  �*  R  R  �*  R  R   '��  �;.  G$  �  �  �*  N$   '��  ��B  G$    &  �*  R  R  N$   '��  ��,  G$  ?  Y  �*  R  R  N$  R     ,!T  q  -�E  �  -�F  �   .�&  .�7  	  �o  >u   �| CG$  /Q  b�   �  /�F c�  /�R  d�  /3  e�  /�  f�  /�K  g�  /�@  h�   0all i�  ?1�� �d  :!  �|*   NF  �+  �E  �n  p0  �+  �%  �+  2S  �+  2�R  �+  23  �+  2�$  �+  2�K  �+  2�@  �+  2�@  �+   �4  �Z  �  �  �*    �=  y)  �  �  �*   3�� �    �*  4+  n   3��   %  �*  N$  n   3�� 5  @  �*  n   3N  P  [  �*  G$   3�� k  v  �*  4+    �  �U  �  �  �*  4+   !�&  �.  2*  �  �  �*    �F  &�;  �  �  �*  :+  �    �9  )�Q  �  �  �*  :+  )+    WR  ,`2      �*  :+  �*    �S  /=  3  C  �*  �*  +   4e  7,  S  �*  +  n    �$  �*   2OD  �*  2gP  �*  2�F  $�*  5< �  6< r�  �  }-  n   7�h  �ܧ  �  48   8�m  �~�  �#  9��  ~�  �#  48    :id ��  �U  �n   2�I  �|*   �  �<?  4  ?  �*  �*   ;id �N  Y  �*  �*   <id �i  o  �*   =4H  ��(  n  �  �*    �o  u�  �  �*   �o  ~�  �  �*  �*   &�o  ��  �  �*  N$   �o  ��  �  �*  �*  N$  �   �o  �  !  �*  �*  �*  �   5  �1  <  �*  G$   *�  ��*  �*  T  _  �*  �*   *H�  ��N  z   w  }  �*   *U  �9  2*  �  �  �*  �*   *2  �t*  2*  �  �  �*  �*   >jP  �D  �  �  �*   8RD  �Q  �*  ?�o  7�  
   �*  �*   @�K  :�N  @�A  =�5  �K  @I  �  <   �    �,  CH<  P   e   �*  �*  �*  �   �  �     �  � >	  <P+  =E+  >[+  @�+  A�+  B,  C+,  DF,  Ef,  F�,  G�,  H�,  �K .!  A�T  1
!  Bok  C'L C�p CFM  D�K !  �-    ד  �R!  ��  �y  � �k  �4  �K*  ,{�  k   E(�  T�  �#  �#   F	L ^�#  Gid  �  HKK Yq  H�L Zq  H�f [&  I&c �!  �!  �,  �,   &&c &�!  �!  �,  n   &&c ,�!  �!  �,  �#  n   J/L 2R!  "  "  �,  G$   K�J 7�K �   R!  >"  g"  -  	-  -  -  -  -  -  !-   �!  K�J FK �   R!  �"  �"  -  	-  -  -  !-   K�L O�L �   R!  �"  �"  -  	-  '-  '-  --  3-  3-  9-   �!  K}I ]cK G$  R!  #  #  -   K<M b�K 2*  R!  :#  @#  -   KK gJ G$  R!  `#  z#  -  	-  '-  '-  n   L�L pxL G$  R!  �#  -    5�I �#  &�J ��#  �#  �-  n   J�J ��#  �#  �#  �-  G$   ,3�  q  ,�e  q  ,�$  &   W�  1�,  R!  Mͳ  � .  N_Tp 7    .   .    O)%  Kk  G$  G$  N$   Pint T$  q  QGT  Pd$  >   �  u$  �  �  o  �	  �  qW  !G$    "�$  �  #  .  <�$  `  DG$  �  W�$  �  _�$  �  eG$  t   mG$  a  uG$    ~G$  �  �G$  3  �G$  �  �G$  H  �G$  y  �G$    �G$  s  �G$  T   �G$  �  �G$  F  �G$  �  �G$  �  �G$    �G$  V  �G$  �  Rs  Nj$  �  Vj$  \	  2G$  o  7G$  �  <G$  �  CG$  �  G$  
&  STpO qO !&  U$   E�)  	�  $,n  -y  K  :�'  �e  =n  � ?k  "  @N$  �4  AK*  �J  BQ*  �A  O�&  �&  W*   �A  Q�&  �&  W*  ]*   �A  V�&  �&  W*  G$   *�
 Y51  V&  �&  �&  c*  n&   *�
 ]�R  b&  '  '  c*  z&   *� c?  V&  0'  @'  W*  J&  &   V_ m.   T'  d'  W*  V&  J&   *�3  q89  J&  |'  �'  c*   V.E  ��3  �'  �'  W*  V&  Q*   V�(  ��(  �'  �'  W*  V&   N_Tp q   >&  WZD  ��)  FF�  �k   H��  �'!  H�4  �=!  H� �2!  %��  �'(  -(  �,   6��  �>(  I(  �,  �,   '*  ��}  �'  b(  h(  �,   'Ư  �?s  	(  �(  �(  �,   '�F  �Ϭ  �,  �(  �(  �,   '�F  ��  �'  �(  �(  �,  G$   'a�  �
�  �,  �(  �(  �,   'a�   ��  �'  )  )  �,  G$   '�:  ,�  �'  &)  1)  �,  �'   '�F  		n  �,  J)  U)  �,  �'   '(*  ��  �'  n)  y)  �,  �'   ' I  h�  �,  �)  �)  �,  �'   '�O  7k  �'  �)  �)  �,  �'   'WC  ]�  �,  �)  �)  �,   ,{�  k  ,�  	   .8E  �'   �� �� �� U2*  7&*  X8�   Y�  Y�  �  �  �  Y	  Yq  YT$  >&  Y�'  �'  �  Y    �   G$  G$    �  	    Y  Y�  Y	  Z7   �*  [ Y    �*  �*  N$  �  Yu   u   �  Ye   e   +  j   k  Z�*  +  [ Z)+  )+  [ /+  �*  Yo   o   7   �l  %   j�  #%   \tm ,,�+  ,g  .G$   �  /G$  �  0G$  ��  1G$  ��  2G$  ��  3G$  ��  4G$  �  5G$  d�  6G$   ��  7%   $~�  8N$  ( Q\�  >P+  Oѯ  H*  ,  E+  E+   O��  ME+  %,  %,   [+  O�  CE+  @,  @,   E+  O#�  ak  [,  [,   a,  [+  O�� fk  {,  {,   �,  E+  O��  W%,  �,  {,   O[v  \%,  �,  {,   O��  R,   �,  k  ,   N$  [,   �'  Y�,  k  �)  Y�'  G$  R!  Y$  $  Y�!  g"  Y-  �!  Y-  �"  Y'-  �!  Y3-  ]Y  M-  W-  ^h  W-   �*  _^�  }-  `w  �G$  `-�  �G$   �  ]�  �-  �-  ^h  �-  a4&  rn   }-  �   b
!  .�-  �-  ^h  �-   �-  �#  ]�#  �-  �-  ^h  �-  `4&  �n   �-  ]�#  .   .  ^h  �-  ^#  �*   Y@+  c$  P.  N_Tp 7   d__a �P.  d__b �U.    .   .  e"  @C   �q.  �.  fh  �.  � g�.  �hDK 8-  �g-  �hWK 9�.  �h"y  :-  �g-  �hL ;�.  � -  	-  -  !-  el"  `C   ��.  2/  fh  �.  � g2/  �h"y  G-  �g-  �hL H7/  � 	-  !-  e�"  pC   �S/  �/  fh  �.  � g�/  �hDK P'-  �g'-  �hWK Q�/  �h"y  R3-  �g3-  �hL R�/  � 	-  --  9-  e�"  �C   ��/  �/  fh  �.  �  e#  �C   ��/  0  fh  �.  �  e@#  �C   �0  v0  fh  �.  � gv0  �hDK h'-  �h�h  i'-  �h�  in  �i�C   j__d kn  �B   	-  ez#  �C   ��0  �0  fh  �.  �  ]�!   �0  �0  ^h  �0  ^#  �*   �,  k�0  �I �CJ   ��0  =1  l�0  � m�-  �C��  3
1  n.  C oD p�-  D   3*1  l.  Sq"D r�C�  r*D:8   k�0  XL 0D   �X1  s1  l�0  � r>D�0  sKDM8   ]�!   �1  �1  ^h  �0  `4&  'n   ks1  8L PDD   ��1  <2  l�1  � l�1  �m�-  RD��  )	2  n�-  HC n�-  gC t�-  RD��  �n�-  HC n�-  gC   p�-  {D   ))2  l.  Sq�D rrD�  r�D:8   ]�!   J2  j2  ^h  �0  `(�  -�#  `4&  -n   k<2  �I �D.   ��2  �2  lJ2  � nS2  �C l^2  �m�-  �D�  /�2  n�-  �C n�-  �C t�-  �D�  �n�-  �C n�-  �C   r�D�   uU  =�2   �$  u�   >�2  uB  ?�2  u�  E%3   �$  uB   F%3  uC  G%3  ue  H%3  u8  I%3  u�  J%3  u

  Xr3   �$  u�  Yr3  u�
  Zr3  v�   `�3  �$  u�  f�3   �$  u�  g�3  u�  h�3  u�  n�3   �$  u�	  o�3  u�  p�3  uH  v�3   �$  u`  w�3  uw  x�3  u   y�3  u~  34   	%  u   �34  u�  �34  u  �34  u�   �34  u�  �34  u�	  �34  u�  ��4   %  u  ��4  u  ��4  u�  ��4  u�  ��4   %  u�  ��4  u�  ��4  u�  ��4  um  ��4   *%  u	  ��4  u2	  ��4  u�  ��4  u9  ��4  u[  �75   5%  uJ  �75  u�  �75  u7  �75  u�  �l5   @%  uI	  �l5  u$	  �l5  u�   ��5   K%  uN  ��5  up  ��5   V%  u�  ��5  u:  ��5  u�  ²5  ud   ò5  u�  ��5   a%  u  ��5  u�  ��5  u�	  �6   l%  u�  �6  u  �96   w%  u�  �96  u�  �96  u�  �96  u+  �n6   �%  u�  �n6  u�   �n6  u  �6   �%  u�
  �6  u�  �6  u  ��6   �%  u   ��6  uF  ��6  u�  ��6   �%  u�  ��6  u�  ��6  uD  O7   �%  u�  P7  u1  Q7  u�  W;7   �%  u^  X;7  u�  3X7   �%  u�  4X7  u�   8u7   �%  u�  9u7  ul	  =�7  �%  uN  >�7  u^  ?�7  uL  @�7  ua  D�7  �%  uB  E�7  u�	  F�7  u  G�7  u  H�7  uy  I�7  u�   8   �%  u�  !8  wx!  �I �EY�#  x>  Y  M8  �%   y�  �1  �%    �3   ��  jM �M �V  ��       (  _� �7   �  �  8k  �{  k   ]�  k  \�   k  �D  !k  �3  "k  U>  #k  &�  $k  �  %k  �*  &k   ڡ  'q  $�U  (q  %TL  )q  &�I  *q  'Q  +q  (�C  ,q  )�J  -q  *1  .k  ,o(  /q  0�U  0q  1PL  1q  2�I  2q  3Q  3q  4�C  4q  5�J  5q  6 q  �  std  �"  5>   6�"  7�"  @t$  	%  0�=  �n  �b  �q  Fe  �"  
�3  �=  �  �(  �(   �  eq �<-  �(    �(  �(   lt ��1  �(  !  �(  �(   ��  eF  �"  E  �(  �(  n   �K  �9  n  _  �(   �(  
!  �(  �  �(  n  �(   1  �A  �(  �  �(  �(  n   �5  �'  �(  �  �(  �(  n   �3  �A  �(  �  �(  n  �   +  :  �  	  �(   �  �C   �P  �  (  �(   �B  $6  �(  G  �(  �(   eof (�:  �  ?  ,N0  �  �(    _� 	�7   �?  	�%   K  
\  �$   �e  
_n  �4  
c�(  �J  
d�(  ��  
q�  �  �(   ��  
s�  �  �(  �(   W  
y�  �(  �"    �  �J  pz  �B  R  �   %  k   �B  A  �(  k  �(    �e  y�  [V  k  R  �G  !   <  x�  �4  {�  �J  |�  �J  5&  `S  �T(  ~J  �z  �J  �  �%  �  �K  �R   I  �R  :!  ��(   %H  ��  �   �3  2k  �G  7�"  t3  B)  �'  ��O  )  V  ��N  �(  [  a  ")   3  �o+  �(  x  ~  ")   �P  ��O  �  �  �(   �M  ��P  �  �  �(   �,  �-  �  �  �(  R   �+  ��R  k  �  �  �(   3  �   k      �(  �(  �(   �/  !�B  �(  6  R  R  �(   �O  �|6  I  T  �(  �(    (  ��6  h  s  �(  �(   !�   �-  k  �  �  �(   "�1  o�*  k  �  �(  �(  R    !�A  $n%  k  �  �  �(   !�A  (�I  k  �  �  �(  k   !"A  ,�%  �(      �(   !�1  2E)  �  -  3  �(   !�/  6;&  �  K  Q  �(    �>  :�>  e  k  �(   !S  A:2  R  �  �  �(  R  �"    �#  K�(  �  �  �(  R  R  �"   !9  S>$  R  �  �  �(  R  R   !-U  [�7  �(  �    �(  �"   #�5  d�-  '  k  �"  R   #	1  m�P  G  k  �"  R   #�3  v\-  g  k  R  q   #nU  ��-  �  k  �  �   #nU  �nG  �  k  �  �   #nU  ��   �  k  k  k   #nU  �IP  �  k  �"  �"   �J  �rR  �"  	  R  R    �=  ��H  	  /	  �(  R  R  R    V  �)  C	  I	  �(   $�'  �D*  )  %�0  �j	  p	  �(   &�0  ��	  �	  �(  �(   �0  ��	  �	  �(  )   �0  ��	  �	  �(  )  R  R   �0  ��	  �	  �(  )  R  R  �(   �0  �
  
  �(  �"  R  �(   �0  �*
  :
  �(  �"  �(   �0  �J
  _
  �(  R  q  �(   %�0  "p
  {
  �(  �"   '�  *,Q  )  �
  �
  �(  )   '�  2�G  )  �
  �
  �(  �"   '�  =�%  )  �
  �
  �(  q   'S� f�&  �       �(   'S� q�>  �    %  �(   (end y<  �  >  D  �(   (end �6;  �  ]  c  �(   'I ��$  �  |  �  �(   'I ��7  �  �  �  �(   '��  �lC  �  �  �  �(   '��  �CM  �  �  �  �(   'r ��R  R  �  �  �(   '�K  �r5  R      �(   '�3  �j=  R  6  <  �(   )�� �  Q  a  �(  R  q   )�� ��F  v  �  �(  R   'I  v  R  �  �  �(   )�E  �|U  �  �  �(  R   )�1  -�  �  �  �(   '�� 5�?  �(  �  �  �(   '�:  D�6  �      �(  R   '�:  UW  �  7  B  �(  R   (at k
/  �  Z  e  �(  R   (at ��7  �  }  �  �(  R   '�F  ��/  )  �  �  �(  )   '�F  �k:  )  �  �  �(  �"   '�F  ��H  )  �  �  �(  q   '@  DA:  )      �(  )   '@  U�1  )  1  F  �(  )  R  R   '@  )�D  )  _  o  �(  �"  R   '@  ��*  )  �  �  �(  �"   '@  �6  )  �  �  �(  R  q   )�G  -aN  �  �  �(  q   *�3  �b*  )  �  �  �(  )   '�3  ^ 2  )    -  �(  )  R  R   '�3  �=  )  F  V  �(  �"  R   '�3  z�T  )  o  z  �(  �"   '�3  � @  )  �  �  �(  R  q   )� ��E  �  �  �(  �  R  q   '� �\+  )  �  �  �(  R  )   '� �u>  )    )  �(  R  )  R  R   '� g|=  )  B  W  �(  R  �"  R   '� "�@  )  p  �  �(  R  �"   '� 9k<  )  �  �  �(  R  R  q   '� K�'  �  �  �  �(  �  q   'bL  d�R  )  �     �(  R  R   'bL  t�2  �    $  �(  �   'bL  �L&  �  =  M  �(  �  �   '�%  �9F  )  f  {  �(  R  R  )   '�%  �|<  )  �  �  �(  R  R  )  R  R   '�%  ��T  )  �  �  �(  R  R  �"  R   '�%  ��A  )  �    �(  R  R  �"   '�%  b>  )  -  G  �(  R  R  R  q   '�%  3%  )  `  u  �(  �  �  )   '�%  'V7  )  �  �  �(  �  �  �"  R   '�%  <�+  )  �  �  �(  �  �  �"   '�%  Q'S  )  �  	  �(  �  �  R  q   '�%  vj.  )  "  <  �(  �  �  k  k   '�%  ��9  )  U  o  �(  �  �  �"  �"   '�%  �C  )  �  �  �(  �  �  �  �   '�%  �>/  )  �  �  �(  �  �  �  �   !�?  ��&  )  �    �(  R  R  R  q   !�1  �O  )    9  �(  R  R  �"  R   ,)  �z-  k  ]  R  q  �(   ++E  �3J  k  �  R  q  �(   '�5  ��)  R  �  �  �(  k  R  R   )n	 @D  �  �  �(  )   'W�  �6  �"  �  �  �(   '�A  %�A  �"      �(   '��  ,Z5  }  %  +  �(   '�(  �;  R  D  Y  �(  �"  R  R   '�(  I�%  R  r  �  �(  )  R   '�(  X�5  R  �  �  �(  �"  R   '�(  �^   R  �  �  �(  q  R   '�(  v�S  R  �  �  �(  )  R   '�(  	K  R    +  �(  �"  R  R   '�(  �o?  R  D  T  �(  �"  R   '�(  J5  R  m  }  �(  q  R   'NW  ��Q  R  �  �  �(  )  R   'NW  /�I  R  �  �  �(  �"  R  R   'NW  ��,  R  �  �  �(  �"  R   'NW  ��;  R    &  �(  q  R   '�S  ��I  R  ?  O  �(  )  R   '�S  >T?  R  h  }  �(  �"  R  R   '�S  05  R  �  �  �(  �"  R   '�S  $S:  R  �  �  �(  q  R   '�>  2hL  R  �  �  �(  )  R   '�>  SUB  R    &  �(  �"  R  R   '�>  Q�2  R  ?  O  �(  �"  R   '�>  _�K  R  h  x  �(  q  R   '�4  qT  R  �  �  �(  )  R   '�4  j�K  R  �  �  �(  �"  R  R   '�4  ��5  R  �  �  �(  �"  R   '�4  N.  R    !  �(  q  R   'U+  �)  	  :  J  �(  R  R   '��  �!1  �"  c  n  �(  )   '��  ��T  �"  �  �  �(  R  R  )   '��  ��O  �"  �  �  �(  R  R  )  R  R   '��  �;.  �"  �  �  �(  �"   '��  ��B  �"    &  �(  R  R  �"   '��  ��,  �"  ?  Y  �(  R  R  �"  R     ,!T  q  -�E  �  -�F  �   .�&  .�7  	  �o  >2   �| C�"  /Q  b�   �  /�F c�  /�R  d�  /3  e�  /�  f�  /�K  g�  /�@  h�   0all i�  ?1�� �d  :!  ��(   NF  �b)  �E  �n  p0  �b)  �%  �n)  2S  �t)  2�R  �t)  23  �t)  2�$  �t)  2�K  �t)  2�@  �t)  2�@  �)   �4  �Z  �  �  ()    �=  y)  �  �  ()   3�� �    ()  �)  n   3��   %  ()  �"  n   3�� 5  @  ()  n   3N  P  [  ()  �"   3�� k  v  ()  �)    �  �U  �  �  ()  �)   !�&  �.  �(  �  �  ()    �F  &�;  �  �  ()  �)  �    �9  )�Q  �  �  ()  �)  �)    WR  ,`2      ()  �)  \)    �S  /=  3  C  ()  \)  h)   4e  7,  S  ()  h)  n    �$  ()   2OD  ()  2gP  ()  2�F  $.)  5< �  6< r�  ]+  n    7id �H  �U  �n   2�I  ��(   �  �<?  �  �  P)  V)   8id �    P)  V)   9id �&  ,  P)   :4H  ��(  n  A  \)    �o  uX  ^  >)   �o  ~n  y  >)  D)   &�o  ��  �  >)  �"   �o  ��  �  >)  D)  �"  �   �o  ��  �  >)  D)  D)  �   5  ��  �  >)  �"   *�  ��*  D)      >)  D)   *H�  ��N  7   4  :  J)   *U  �9  �(  R  ]  J)  D)   *2  �t*  �(  u  �  J)  D)   ;jP  �D  �  �  D)   <RD  �Q  D)  =�o  7�  �  >)  ()   >�K  :�N  >�A  =�5  �K  @I  �  �  �    �,  CH<     "   >)  D)  D)  �   �  �     �  � >	  <�)  =�)  >�)  @G*  AR*  Bl*  C�*  D�*  E�*  F�*  G�*  H+  ?�  H!  @Sv  L�   �O  L0+    AQ�   B��   B+�  B�1   �  N�   �   ��  Y�"  CFv  ^��  �   q  q  q    ד  �T!  ��  �y  � �k  �4  ��(  ,{�  k   D��  �!  3ҽ  zm!  x!  �+  n   ,!T  q  E�  �(   5�  �!  F�q  -Y�  �!  �!  �+  �!  �"   Ge�  `�!  �!  �!  �+  �"   ,!T  q  E�  �(   W�  1�+  D
�  0"  3ҽ  z"  "  �,  n   ,!T  q  E�  �(    H��  F�q  G��  I"  Y"  �,  �!  �"   Ge�  d0"  n"  y"  �,  �"   ,!T  q  E�  �(     I)%  Kk  �"  �"  �"   Jint �"  q  KGT  P�"  >   �  �"  �  �  o  �	  �  qW  !�"    "#  �  #  .  <�"  `  D�"  �  W�"  �  _#  �  e�"  t   m�"  a  u�"    ~�"  �  ��"  3  ��"  �  ��"  H  ��"  y  ��"    ��"  s  ��"  T   Ȩ"  �  Ш"  F  ר"  �  �"  �  �"    �"  V  �"  �  Ls  N�"  �  V�"  \	  2�"  o  7�"  �  <�"  �  C�"  �  �"  k$  MNpO qO !l$  O$   E_(  	�  $,n  -y  K  :0&  �e  =n  � ?k  "  @�"  �4  A�(  �J  B�(  �A  O�$  �$  �(   �A  Q%  %  �(  �(   �A  V(%  3%  �(  �"   *�
 Y51  �$  K%  V%  �(  �$   *�
 ]�R  �$  n%  y%  �(  �$   *� c?  �$  �%  �%  �(  �$  e$   F_ m.   �%  �%  �(  �$  �$   *�3  q89  �$  �%  �%  �(   F.E  ��3  �%  &  �(  �$  �(   F�(  ��(  &  &&  �(  �$   P_Tp q   �$  ?ZD  �T(  QF�  �k   R��  �)!  R�4  �?!  R� �4!  %��  ��&  �&  @+   S��  ��&  �&  @+  F+   '*  ��}  ]&  �&  �&  Q+   'Ư  �?s  j&  �&  �&  Q+   '�F  �Ϭ  W+  '  '  @+   '�F  ��  5&   '  +'  @+  �"   'a�  �
�  W+  D'  J'  @+   'a�   ��  5&  c'  n'  @+  �"   '�:  ,�  ]&  �'  �'  Q+  P&   '�F  		n  W+  �'  �'  @+  P&   '(*  ��  5&  �'  �'  Q+  P&   ' I  h�  W+  �'  �'  @+  P&   '�O  7k  5&  (  "(  Q+  P&   'WC  ]�  F+  ;(  A(  Q+   ,{�  k  ,�  	   .8E  5&   �� �� �� O2*  7�(  T8�   U�  U�  �  �  �  U	  Uq  U�"  �$  U0&  0&  �  U    �   �"  �"    �  	    U  U�  U	  V7   ")  W Y    3)  9)  �"  �  U2   2   �  U"   "   h)  '   k  V\)  )  W V�)  �)  W �)  \)  U,   ,   �l  %   j�  #%   Xtm ,,G*  ,g  .�"   �  /�"  �  0�"  ��  1�"  ��  2�"  ��  3�"  ��  4�"  �  5�"  d�  6�"   ��  7%   $~�  8�"  ( K\�  >�)  Iѯ  Hf(  l*  �)  �)   I��  M�)  �*  �*   �)  I�  C�)  �*  �*   �)  I#�  ak  �*  �*   �*  �)  I�� fk  �*  �*   �*  �)  I��  W�*  �*  �*   I[v  \�*  +  �*   I��  R,   0+  k  ,   �"  �*   Vq  @+  Y$   5&  UL+  k  Y(  U5&  �  Z�  q+  �+  [h  �+  \4&  rn   ]+  ]�   (�D   ��+  ^q  �^q  �^q  � T!  Z]!  �+  �+  [h  �+  \4&  zn   �+  �!  �"  _�!  �D*  �,  �,  `h  �,  � ^�!  �^�"  �aVE   E,  b__i An  �C  c�+  �E|   1�,  d�+   e�+  Pfc+  �E   �dz+   eq+  P  g�E�3   �+  �!  Z"  �,  �,  [h  �,  \4&  zn   �,  0"  _5"  F*  ��,  a-  `h  a-  � ^�!  �^�"  �a�F   -  b__i [n  D  c�,  �F|   KW-  d�,   e�,  Pfc+  �F   �dz+   eq+  P  g�F�3   �,  Z�!   t-  �-  [h  �,  [#  �(   hf-  /N @GB   ��-  �-  et-  � ioGjzGg�G�3   kf-  MM �G   ��-  �-  et-  � g�G�-  l�G�3   ZY"   .  .  [h  a-  [#  �(   h�-  N �GB   �0.  L.  e.  � i�Gj�Gg�G�3   k�-  LN  H   �g.  �.  e.  � gH.  lH�3   mU  =�.   #  m�   >�.  mB  ?�.  m�  E�.   (#  mB   F�.  mC  G�.  me  H�.  m8  I�.  m�  J�.  m

  X/   3#  m�  Y/  m�
  Z/  n�   `-/  >#  m�  f>/   I#  m�  g>/  m�  h>/  m�  ng/   T#  m�	  og/  m�  pg/  mH  v�/   _#  m`  w�/  mw  x�/  m   y�/  m~  �/   j#  m   ��/  m�  ��/  m  ��/  m�   ��/  m�  ��/  m�	  ��/  m�  �0   u#  m  �0  m  �0  m�  �0  m�  �S0   �#  m�  �S0  m�  �S0  m�  �S0  mm  ��0   �#  m	  ��0  m2	  ��0  m�  ��0  m9  ��0  m[  ��0   �#  mJ  ��0  m�  ��0  m7  ��0  m�  ��0   �#  mI	  ��0  m$	  ��0  m�   �'1   �#  mN  �'1  mp  �D1   �#  m�  �D1  m:  �D1  m�  �D1  md   �D1  m�  Ʌ1   �#  m  ʅ1  m�  ˅1  m�	  Ѯ1   �#  m�  Ү1  m  ��1   �#  m�  ��1  m�  ��1  m�  ��1  m+  � 2   �#  m�  � 2  m�   � 2  m  �)2   �#  m�
  �)2  m�  �)2  m  �R2   �#  m   �R2  mF  �R2  m�  �{2   $  m�  �{2  m�  �{2  mD  O�2   $  m�  P�2  m1  Q�2  m�  W�2   #$  m^  X�2  m�  3�2   .$  m�  4�2  m�   83   9$  m�  93  ml	  =$3  D$  mN  >$3  m^  ?$3  mL  @$3  ma  DY3  O$  mB  EY3  m�	  FY3  m  GY3  m  HY3  my  IY3  m�   �3   Z$  m�  !�3  +�  ��  $  �3  n   o>  Y  �3  $   p�  �1  $    �   v�  [R 	f �b ��       (  _� �7   �  #  �� �  �  �  c   �  �  u   �  �O �   o  �O �   �	  pW   �   �  qW  !�   int   "�   �    #>   ` &u   ` 'c   �^ (�   �^ )�   �T *�   �T +�   iY ,>   hY -�   �e 0u   �e 1c   [ 2�   [ 3�   Q 4�   Q 5�   �_ 6>   �_ 7�   �] :�   �] ;�   �Q >>   �Q ?�   Fd �   .  <�   `  D�   �  W�   �  _�   �  e�   t   m�   a  u�     ~�   �  ��   3  ��   �  ��   H  ��   y  ��     ��   s  ��   T   Ƚ   �  н   F  ׽   �  �   �  �     �   V  �   Q   �  s  NX   �  VX   \	  2�   o  7�   �  <�   �  C�   �  �   X   	\  �   gX  �   X\  &<  	X\  X,Q  
$Z  .�   
\ /X   
� 1  
Z  2,   
K]  3X   
�_  4,   
\W  5,   
�Z  6,   
-_  8p   
VY  9�  $
`  :�  (
�Y  ;�  ,
7_  <�  0
BY  =	  4
b\  >�  8
\  ?�  <
7Y  @�  @
 Z  A  D
SX  B  H
n4 D�   L
`  Fj  P
*5 Gj  T &  j  �  ,   j   <  Q  &  �  �  ,   j   �  v  �   �  j    �    �    �  j   �  �   �  j   �  j  �  �  �  j     Q   �    j     pO qO !   std . SC  @(  v  6�  x  K�  
�  M�   x  Ow  �  SC  �   �  Qw  �  �  SC   �  R  �  �  SC     T8  �  �  �  YC   x  Z�  �  SC   x  \�    SC  _C   x  _    SC  �   x  c-  8  SC  eC   �  p�  kC  P  [  SC  _C   �  t�  kC  s  ~  SC  eC   �  {�  �  SC  �    n	 ~%  �  �  SC  kC   �  ��  qC  �  �  YC   �  �h  xC  �  YC    P   :P  �  �L   � 	  �S 0L %  '0	�=  �	  �b  �Q   Fe  �   �#  �	  �&  �
  �f �(  !�3  �=    'E  -E   .  "eq �<-  qC  �  -E  -E   "lt ��1  qC  �  -E  -E   #��  eF  �   �  3E  3E  �
   #�K  �9  �
  �  3E   #�(  
!  3E     3E  �
  -E   #1  �A  9E  D  9E  3E  �
   #�5  �'  9E  h  9E  3E  �
   #�3  �A  9E  �  9E  �
  .   #+  :  .  �  ?E   9  #�C   �P  9  �  -E   #�B  $6  qC  �  ?E  ?E   $eof (�:  9  %?  ,N0  9  ?E    E  �	  9Q  p
  
G0  s
   
�T  t(  %  {J	  P	  �J   %  �`	  k	  �J  
   �:  �b;  
  �	  �	  �J   �T  �4>  �	  �	  �J  (   �T  �QM  (  �	  �	  �J   �F  ��?  �J  �	  �	  �J  
    I  �O  �J  
  
  �J  
   (*  �	H  	  $
  /
  �J  
   �O  �eT  	  G
  R
  �J  
   �O  ́?  
  j
  u
  �J  �J   &�$  (   �:  Z>   _� �7   0j   1�   2�   3�   59  6O  7e  8{  :�   ;�   <  =#  ?�  @�  BX   C|   D�   E�   GD  HZ  Ip  J�  L�   M  N  O.  Q�  R�  5SE  6�F  7�F  �?  �%   K  \�  '�C   (�e  _�
  (�4  c�F  (�J  d�F  ��  q�  �  �F   ��  s�  �  �F  �F   )W  y�  �F  �     y  �J  p%  *�B  G  +y   ,%  �   -�B  6  �F  �  �F    (�e  y�  .[V  `  G  ,�G  !
   (<  xy  (�4  {�  (�J  |�  (�J  �D  (`S  ��D  (~J  �%  (�J  �#%  	�%  ��  
�K  �G   
I  �G  
:!  ��F   	%H  ��  +�   /�3  2`  /�G  7  /t3  B-G  0�'  ��O  G  V  ��N  qC  P  V  8G   3  �o+  qC  m  s  8G   �P  ��O  �  �  G   �M  ��P  �  �  G   �,  �-  �  �  G  G   �+  ��R  �  �  �  G   3  �   �  �    G  �F  �F   #�/  !�B  G  +  G  G  �F   �O  �|6  >  I  G  �F   1(  ��6  ]  h  G  �F   2�   �-  �  �  �  G   3�1  o�*  �  �  G  �F  G    2�A  $n%  �  �  �  G   2�A  (�I  �  �  �  	G  �   2"A  ,�%  G    
  G   2�1  2E)  �  "  (  G   2�/  6;&  �  @  F  G   1�>  :�>  Z  `  	G   2S  A:2  G  x  �  G  G  �   1�#  K�(  �  �  G  G  G  �   29  S>$  G  �  �  G  G  G   2-U  [�7  qC  �  �  G  �   4�5  d�-    �  �  G   4	1  m�P  <  �  �  G   4�3  v\-  \  �  G  Q    4nU  ��-  |  �  �  �   4nU  �nG  �  �  �  �   4nU  ��   �  �  �  �   4nU  �IP  �  �  �  �   #�J  �rR  �   �  G  G   1�=  ��H    $  	G  G  G  G   1V  �)  8  >  	G   5�'  �D*  G  6�0  �_  e  	G   7�0  �v  �  	G  �F   6�0  ��  �  	G  G   6�0  ��  �  	G  G  G  G   6�0  ��  �  	G  G  G  G  �F   6�0  ��    	G  �  G  �F   6�0  �%  5  	G  �  �F   6�0  �F  [  	G  G  Q   �F   6�0   l  w  	G  !G   6�0  �  �  	G  -%  �F   6�0  "�  �  	G  �    8�  *,Q  'G  �  �  	G  G   8�  2�G  'G  �  �  	G  �   8�  =�%  'G       	G  Q    8�  Mo_ 'G  9  D  	G  !G   8�  Y.c 'G  ]  h  	G  -%   8S� f�&  �  �  �  	G   8S� q�>  �  �  �  G   9end y<  �  �  �  	G   9end �6;  �  �  �  G   8I ��$  �  �    	G   8I ��7  �    "  G   8��  �lC  �  ;  A  	G   8��  �CM  �  Z  `  G   8)^ �^\ �  y    G   8%] ��a �  �  �  G   8hf �*] �  �  �  G   8wY �Je �  �  �  G   8r ��R  G  �  �  G   8�K  �r5  G      G   8�3  �j=  G  3  9  G   :�� ��  N  ^  	G  G  Q    :�� ��F  s  ~  	G  G   :be  VT �  �  	G   8I  v  G  �  �  G   :�E  &|U  �  �  	G  G   :�1  -�  �  �  	G   8�� 5�?  qC      G   8�:  D�6  �  +  6  G  G   8�:  UW  ~  O  Z  	G  G   9at k
/  �  r  }  G  G   9at ��7  ~  �  �  	G  G   8��  ��O ~  �  �  	G   8��  �}Y �  �  �  G   8�G  �@\ ~  �  �  	G   8�G  �e �      G   8�F  ��/  'G  5  @  	G  G   8�F  �k:  'G  Y  d  	G  �   8�F  ��H  'G  }  �  	G  Q    8�F  �x` 'G  �  �  	G  -%   8@  �A:  'G  �  �  	G  G   8@  ��1  'G  �  �  	G  G  G  G   8@  ��D  'G    '  	G  �  G   8@  ��*  'G  @  K  	G  �   8@  �6  'G  d  t  	G  G  Q    8@  �] 'G  �  �  	G  -%   :�G  -aN  �  �  	G  Q    8�3  <b*  'G  �  �  	G  G   8�3  Ipf 'G  �     	G  !G   8�3  ^ 2  'G    .  	G  G  G  G   8�3  n�=  'G  G  W  	G  �  G   8�3  z�T  'G  p  {  	G  �   8�3  � @  'G  �  �  	G  G  Q    8�3  ��a 'G  �  �  	G  -%   :� ��E  �  �  	G  �  G  Q    :� ��V     	G  �  -%   8� �\+  'G  0  @  	G  G  G   8� �u>  'G  Y  s  	G  G  G  G  G   8� |=  'G  �  �  	G  G  �  G   8� "�@  'G  �  �  	G  G  �   8� 9k<  'G  �  �  	G  G  G  Q    8� K�'  �    !  	G  �  Q    8bL  d�R  'G  :  J  	G  G  G   8bL  t�2  �  c  n  	G  �   8bL  �L&  �  �  �  	G  �  �   :H�  �M\ �  �  	G   8�%  �9F  'G  �  �  	G  G  G  G   8�%  �|<  'G  �    	G  G  G  G  G  G   8�%  ��T  'G  1  K  	G  G  G  �  G   8�%  ��A  'G  d  y  	G  G  G  �   8�%  b>  'G  �  �  	G  G  G  G  Q    8�%  3%  'G  �  �  	G  �  �  G   8�%  'V7  'G  �    	G  �  �  �  G   8�%  <�+  'G  &  ;  	G  �  �  �   8�%  Q'S  'G  T  n  	G  �  �  G  Q    8�%  vj.  'G  �  �  	G  �  �  �  �   8�%  ��9  'G  �  �  	G  �  �  �  �   8�%  �C  'G  �    	G  �  �  �  �   8�%  �>/  'G     :  	G  �  �  �  �   8�%  �b 'G  S  h  	G  �  �  -%   2�?  ��&  'G  �  �  	G  G  G  G  Q    2�1  �O  'G  �  �  	G  G  G  �  G   #,)  �z-  �  �  G  Q   �F   #+E  �3J  �    G  Q   �F   8�5  �)  G  -  B  G  �  G  G   :n	 @D  W  b  	G  'G   8W�  �6  �  {  �  G   8�A  %�A  �  �  �  G   8��  ,Z5  r  �  �  G   8�(  <;  G  �  �  G  �  G  G   8�(  I�%  G        G  G  G   8�(  X�5  G  /   ?   G  �  G   8�(  i^   G  X   h   G  Q   G   8�(  v�S  G  �   �   G  G  G   8�(  �K  G  �   �   G  �  G  G   8�(  �o?  G  �   �   G  �  G   8�(  �J5  G  !  !  G  Q   G   8NW  ��Q  G  *!  :!  G  G  G   8NW  ��I  G  S!  h!  G  �  G  G   8NW  ��,  G  �!  �!  G  �  G   8NW  ��;  G  �!  �!  G  Q   G   8�S  ��I  G  �!  �!  G  G  G   8�S  T?  G  �!  "  G  �  G  G   8�S  05  G  *"  :"  G  �  G   8�S  $S:  G  S"  c"  G  Q   G   8�>  2hL  G  |"  �"  G  G  G   8�>  CUB  G  �"  �"  G  �  G  G   8�>  Q�2  G  �"  �"  G  �  G   8�>  b�K  G  �"  #  G  Q   G   8�4  qT  G  %#  5#  G  G  G   8�4  ��K  G  N#  c#  G  �  G  G   8�4  ��5  G  |#  �#  G  �  G   8�4  �N.  G  �#  �#  G  Q   G   8U+  �)  �  �#  �#  G  G  G   8��  �!1  �   �#  $  G  G   8��  ��T  �   $  0$  G  G  G  G   8��  ��O  �   I$  h$  G  G  G  G  G  G   8��  	;.  �   �$  �$  G  �   8��  (	�B  �   �$  �$  G  G  G  �   8��  C	�,  �   �$  �$  G  G  G  �  G   �  &!T  Q   ;�E  "  ;�F  y   %  � >�  �&  �7  �  Qf �o  >�*  (�| C�   <Q  bW%   >%  <�F cW%  <�R  dW%  <3  eW%  <�  fW%  <�K  gW%  <�@  hW%   =all iW%  ?>�� �(  ,:!  ��F   ,NF  �xG  ,�E  ��
  ,p0  �xG  ,�%  ��G  ?S  ��G  ?�R  ��G  ?3  ��G  ?�$  ��G  ?�K  ��G  ?�@  ��G  ?�@  ��G  1�4  �Z  n&  t&  >G   1�=  y)  �&  �&  >G   @�� �&  �&  >G  �G  �
   @�� �&  �&  >G  �  �
   @�� �&  �&  >G  �
   @N  �&  '  >G  �    @�� '  '  >G  �G   1�  �U  3'  >'  >G  �G   2�&  �.  qC  V'  \'  >G   1�F  &�;  p'  �'  >G  �G  >%   1�9  )�Q  �'  �'  >G  �G  �G   1WR  ,`2  �'  �'  >G  �G  rG   1�S  /=  �'  �'  >G  rG  ~G   Ae  7,  �'  >G  ~G  �
    ,�$  >G   ?OD  >G  ?gP  >G  ?�F  $DG  < Bid ��(  ,�U  ��
   ?�I  ��F  1�  �<?  }(  �(  fG  lG   Cid ��(  �(  fG  lG   Did ��(  �(  fG   E4H  ��(  �
  �(  rG    �o  u�(  �(  TG   �o  ~�(  )  TG  ZG   F�o  �)   )  TG  �   �o  �0)  E)  TG  ZG  �  >%   �o  �U)  j)  TG  ZG  ZG  >%   5  �z)  �)  TG  �    �  ��*  ZG  �)  �)  TG  ZG   H�  ��N  %  �)  �)  `G   U  �9  qC  �)  �)  `G  ZG   2  �t*  qC  *  *  `G  ZG   GjP  �D  2%  '*  ZG   HRD  �Q  ZG  I�o  7H*  S*  TG  >G   J�K  :�N  J�A  =�5  #�K  @I  >%  �*  >%   1�,  CH<  �*  �*  TG  ZG  ZG  >%   C(  >(  �%   2%  KW  3R+  L�4  L�$  Lq-  Lc=  Lo'  L�5   L�%  � L�8  �LX)  �L�%  �L�  �LaO  �LY=  � LP  �� L�C  ��LwS  �L�O  � L�?  �L�5  �� K
$ g�+  L)W  L�   L�U  L�A  L�8  L�P   LEH  �� K�4  ��+  LO   L�7  L(  L�Q  LG  �� K��  ��+  L�R   L�-  L�1  LlO  �� Mb4 �-  N�9  iR+  N�N  ��+  N�  J�+  (�P  ��*  O�4  ),  ,  Pdec ),  Ot-  ),  Phex ),  Or'  ),  O< ),   Poct ),  @O� ),  �Q[)  ),   Q�%  "),   Q�  &),   QdO  )),   Q\=  ,),   Q�P  /),    Q�C  3),   @OzS  6),  �O�O  9),  JQ�?  <),  O�7  N2-  ,  O(  Q2-  O�Q  V2-  OO  Y2-   Papp lo-  �+  Pate oo-  Pin wo-  Pout zo-  O�P  }o-   Pbeg ��-   �+  Pcur ��-  Pend ��-   M�8  n.  6�  
��-  .  \L  �   �J   F�  
T.  *.  \L  �   �J  �L   ({'  
E/  R�@  
]�-  K.  [.  \L  �   �J   &!T  Q   ;�E  "   M�Y  /  R�% 	gn.  �.  �.  �L  �   �J   6̾ 	^�.  �.  �L  �   �J   F̾ 	]�.  �.  �L  �   �J  5�   ({'  	E/  &!T  Q   ;�E  "   M�M  
1  8�* �_e  �J  #/  )/  �J   (�b  �Q   8�* �e  �J  N/  T/  �J   8% ��" �J  m/  s/  �J   :cb  �Pc  �/  �/  QK  �    8�-  P  �J  �/  �/  �J   8� � �J  �/  �/  �J   :� !4  �/  �/  QK  �    8�-  �  �J  
0  0  �J   RZ  �/  %0  00  QK  �    :��  �R�  E0  Z0  QK  �J  �J  �J   6�B �k0  q0  QK   :��  +�  �0  �0  QK  �J  �J   &!T  Q   ;�E  "  S�W  "O`@ H4  /  �0  �0  QK  J�  H4   )/  T�W  "-�A H4  /  �0  QK  �J  H4    �K .81  U�T  1Vok  L'L L�p LFM   b1  c�G  e�G  f�G  g�G  h
H  i H  j5H  kKH  llH  m�H  q�H  r�H  t�H  u
I  v0I  xFI  y\I  |hI  ~}I  ��I  ��I  ��I  ��I  ��I  �
J  �J  �*J  �   5-4  
  8EJ   
��   ;qC  �  >02  ;2  KJ  QJ   @�   Ad�  KJ  S2  h2  KJ  �  �+  �    &�   Dx�  KJ  �2  �2  KJ  EJ  �+   &�   G( KJ  �2  �2  KJ  �   �+   <_   JG�  KJ  �2  �2  KJ   �   M��  qC  �2  �2  WJ   Wfd  P� �   3  3  KJ   QY   S� EJ  )3  /3  KJ   �  U?3  J3  KJ  �    �W   X" H4  b3  r3  KJ  �  H4   f  [� H4  �3  �3  KJ  �  H4  �  H4   �W   _: H4  �3  �3  KJ  �  H4   09   b��  
  �3  �3  KJ  
  �+   �  e  �   4  4  KJ   ��   h��  H4  &4  KJ    �^  !-1  � !*�F  �1  �>  bn  X��  `H/  �9  '/   Y\ ]84   (�c T�1  YNY  `w4  $Y�% c�+  ,(�f UZ  Y�b f�4  0Y�R k�4  1YQX o�4  2(�b  LQ   YU r]J  4Y�W y�
  8Y�V |qC  <Y�V �qC  =Y�] �qC  >Y{O ��4  ?Y�Q �]J  @Y9_ �]J  DY�S �qC  H(Q] V�9  Y#c �cJ  LQ5  Y�Z ��  PY�S �H4  TY�T ��  XY�] ��  \(Fe  N9  (�#  OD  (�&  PO  ({'  R/  (��  SS4  ue ��S �5  �5  iJ   ^_ \ 6  6  iJ   �	 N#6  )6  iJ   R�	 �S4  >6  I6  iJ  �    �  ���  qC  a6  g6  oJ   @�  ]�^ uJ  6  �6  iJ  �  �+   8@�  �O uJ  �6  �6  iJ  �F  �+   <_  ��  uJ  �6  �6  iJ   Y /& �6  �6  iJ   �X =�Y 7  
7  iJ   S��  �+[ H4  S4  *7  07  iJ   S�[  ��[ �5  	S4  P7  V7  iJ   ZZ  j` �5  S4  w7  �7  iJ  �5   ZP� �_ �5  S4  �7  �7  iJ  �5   8Tg �oc qC  �7  �7  iJ  �  H4   ZY@ ��e {J  S4  �7  8  iJ  ]J  H4   Z09  ��Q �5  S4  )8  >8  iJ  �5  �+  �+   Z=H  mT �5  S4  _8  o8  iJ  �5  �+   8SR U �5  �8  �8  iJ  �5  �+  �4   8Wc .5O �   �8  �8  iJ  �J   Z� ~ X �   S4  �8  �8  iJ   [�= �iN S4  9  9  iJ  ZG   Z�W  %MZ H4  S4  19  A9  iJ  �  H4   Z�W  }�a H4  S4  b9  r9  iJ  �  H4   8{_ AR qC  �9  �9  iJ   : �< �9  �9  iJ  H4   �5  �4  &!T  Q   ;�E  "   (�  S4  \a ��n.  |;  'n.   N��  �S4  ,�_ ��9  61^ �:  +:  �J  �   �J   71^ �<:  V:  �J  �   �J  �  �+   71^ �g:  �:  �J  �   �J  �F  �+   ]0^ ��9  �:  �:  �J  �   �J   83F   gX �J  �:  �:  �J   8�  yP qC  �:  �:  �J   8�  d qC  �:  ;  �J   :@�  �` ;  );  �J  �  �+   :@�  1�P >;  N;  �J  �F  �+   :<_  C;S c;  i;  �J   &!T  Q   ;�E  "   �9  \�V �Z�-  %=  '�-   N��  eS4  ,�_ i�;  6�a t�;  �;  �J  �   �J   7�a ��;  �;  �J  �   �J  �  �+   7�a �<  *<  �J  �   �J  �F  �+   ]�a ��;  @<  P<  �J  �   �J   83F  �4Y �J  i<  o<  �J   8�  �a[ qC  �<  �<  �J   8�  �5W qC  �<  �<  �J   :@�  �4P �<  �<  �J  �  �+   :@�  �Z �<  �<  �J  �F  �+   :<_  ��Y =  =  �J   &!T  Q   ;�E  "   �;  \gd �n.  �>  '�>   N��  S4  ,�_ B=  6^ &m=  }=  �J  �   �J   7^ 3�=  �=  �J  �   �J  �  �+   7^ B�=  �=  �J  �   �J  �F  �+   ]^ Q*=  �=  �=  �J  �   �J   83F  \�Z �J  >  >  �J   8�  de qC  1>  7>  �J   8�  jkW qC  P>  V>  �J   :@�  y�U k>  {>  �J  �  �+   :@�  ��W �>  �>  �J  �F  �+   :<_  �YQ �>  �>  �J   &!T  Q   ;�E  "   M$ W?  6l* 	>�>  �>  ׀  �   �J   7l* 	4	?  ?  ׀  �   �J  QK   ]k* 	;�>  4?  D?  ׀  �   �J   &!T  Q   ;�E  "   M�E  "@  �M  ��B  ,  x?  ~?  �K   ]`V  W?  �?  �?  0L  �    6aV  ��?  �?  0L   eU  ��4  �?  �?  0L  ,   &!T  Q   ;�E  "  i3 #~P4  �?  @  0L  QK   ^�1  #)�%  @  0L  ,    *=  	  /  W?  _�*  ��+  P@  �+  �+   _*  sR+  j@  R+  R+   _�] .*O  �@  &�R  �9  0O   �9  M�I +B  �� � Q �   �@  �@  UO   �L ۛX �   �@  �@  UO   ?M ��Z qC  �@  �@  UO   Win ĒU 0A  A  0A  UO  �O  �O  �O  �O  �O  �O  �O   (�T  I1  (�f L(  MA  (�L KQ   (KK JQ   Wout t�\ 0A  }A  �A  UO  �O  �P  �P  �P  �P  �P  �P   YA  �K  ��f �   �A  �A  UO  �O  �O  �O  �
   �J ��_ 0A  �A  B  UO  �O  �P  �P  �P   &3�  Q   &�e  Q   &�$  (   �@  _ͳ  �iP  SB  `_Tp 7   iP  iP   _�*  wR+  mB  R+  R+   _;] �qC  �B  &�$  (  �J  �J   _�b  R  �B  `_Tp %   �R  �R   _�   �qC  �B  &�$  (  �J  �J   H4  �
  a	[ 0O�B     b	@  $8�N  !t4 $_�/ C  �   cα  %h/�  qC  4C  &�R  �9  ZG   d�  %��u  *O  &�R  �9  ZG    P  �  e�  fP  eP  �    $   &��D   �  ($),�
  )-n  K  ):�D  (�e  )=�
  (� )?�  ("  )@�  (�4  )A�F  (�J  )B�F  �A  )O�C  �C  �F   �A  )QD  D  �F  �F   �A  )V'D  2D  �F  �    �
 )Y51  �C  JD  UD  �F  �C   �
 )]�R  �C  mD  xD  �F  �C   � )c?  �C  �D  �D  �F  �C  �   _ )m.   �D  �D  �F  �C  �C   �3  )q89  �C  �D  �D  �F   `_Tp Q    �C  ZD  8E   �� �� qC  7   2*  '7'E  g'8   e.  e    .  e�  Ye �[ 	�  8*�F  
�{  *�   
]�  *�  
\�  * �  
�D  *!�  
�3  *"�  
U>  *#�  
&�  *$�  
�  *%�  
�*  *&�   
ڡ  *'Q   $
�U  *(Q   %
TL  *)Q   &
�I  **Q   '
Q  *+Q   (
�C  *,Q   )
�J  *-Q   *
1  *.�  ,
o(  */Q   0
�U  *0Q   1
PL  *1Q   2
�I  *2Q   3
Q  *3Q   4
�C  *4Q   5
�J  *5Q   6 _)%  *K�  �F  �   �   hGT  *P�F  SE  ��  +!�   �  , �   eQ   e  �C  e�D  �D  y  e�    �   e%  
  (%  �  �  e�  e(%  f�  e�  i7   8G  j �$  �%  IG  OG  �  2%  e�*  �*  C(  e�*  �*  ~G  �*  �  irG  �G  j i�G  �G  j �G  rG  e�*  �*  %   �^  -!  kZ  -1�G  �G   1  _aY  -��   �G  �G   l\  -C�   
H  �G   lxZ  -M�    H  �G   _`  -��   5H  �G   l�^  -r�   KH  �G   l_X  -��   fH  �G  fH   �G  l�_  -��  �H  �  �   �G   _�\  -��G  �H  �  �   l4Z  -�,   �H  �  ,   ,   �G   _7`  -��G  �H  �  �  �G   l>]  -	�   
I  �G  %   �    l�Z  -�   %I  �G  %I   +I  �G  l�Y  - %   FI  �G   l�Y  -��   \I  �G   m\  -��   _�_  0�  }I  �   k�]  -W�I  �   _D[  -T�   �I  �   _�[  -a�   �I  �  �   k�\  -)�I  �G   nY@ -��I  �G  �   _�[  -½   
J  �G  �  �   ,    h�]  -i�G  _D]  -w�  *J  �   l}W  -��   EJ  �   �G   -4  �1  84  C4  �4  j5  S4  �9  �5  �5  e�4  �9  �  �9  |;  �;  �;  %=  *=  B=  "@  	  '@  e	  e'@  )/  ,@  o
/  �J  �J  ph  �J   �J  o5/  K  K  ph  �J   oT/  *K  4K  ph  �J   o�  BK  LK  ph  LK   G  /  os/  eK  {K  ph  {K  q__n ��    QK  o�/  �K  �K  ph  �J   o�/  �K  �K  ph  �J   o�/  �K  �K  ph  {K  q__n !�    o�/  �K  �K  ph  �J   1@  o`?   L  
L  ph  
L   �K  o0  L  0L  ph  {K  p#  �F   W?  o~?  DL  WL  ph  WL  p#  �F   0L  �-  o�-  pL  �L  ph  �L  p#  �F  p�!  �L   \L  �J  n.  ow.  �L  �L  ph  �L  p#  �F  p�!  �L   �L  �J  *.  o.  �L  M  ph  �L  p#  �F  p�!  M  r(  
T�L   �J  o6.  M  :M  ph  �L  p#  �F  p�!  :M   �J  s�  VM  q__c VM   ?E  s�  rM  q__c  rM   -E  s�  �M  thR  $�M  tmR  $�M   ?E  ?E  u�  o�8  �M  �M  ph  �M  vw�&  ��   vwY�  ��9     iJ  s�  �M  q__c ,�M   ?E  s6@   N  x__a ��+  x__b ��+   o00  .N  \N  ph  {K  t�  ��J  t;�  ��J  tP�  ��J   o�5  jN  tN  ph  �M   o�5  �N  �N  ph  �M   oZ0  �N  �N  ph  {K   oI6  �N  �N  ph  �N   oJ  o�6  �N  �N  ph  �M   sP@  �N  x__a sR+  x__b sR+   oq0  O  *O  ph  {K  tM�  +�J  tu�  +�J   e�@  �@  sj@  UO  &�R  �9  x__f .0O   +B  o�@  iO  sO  ph  sO   UO  o�@  �O  �O  ph  sO   o�@  �O  �O  ph  sO   sD  �O  t�e  9E  t�e  3E  q__n �
   e<A  HA  e�O  YA  e�O  o�@  P  ZP  ph  sO  r�%  �ZP  rDK ��O  r�Q ��O  rWK �_P  r"y  ��O  rfc ��O  rL �dP   �O  �O  �O  eE  s0B  �P  `_Tp 7   x__a P  x__b P   iP  iP  �A  e�P  MA  e�P  oeA  �P   Q  ph  sO  r�%  t Q  rDK t�P  r�Q u�P  rWK u%Q  r"y  v�P  rfc v�P  rL w*Q   �O  �P  �P  o�	  =Q  RQ  ph  RQ  r�S �(   �J  ok	  eQ  oQ  ph  oQ   �J  oP	  �Q  �Q  ph  RQ  rQ  �
   sSB  �Q  x__a wR+  x__b wR+   smB  �Q  &�$  (  r\C  ��Q  r?)  ��Q   �J  �J  o�	  �Q  R  ph  oQ   o�A  R  HR  ph  sO  r�%  �HR  rDK ��O  r�h  ��O  r�  ׊
   �O  o�8  [R  R  ph  �M  t�%  /R  vw�d 8�F    �J  e�G  s�B  �R  `_Tp %   x__a ´R  x__b ¹R   �R  �R  o�A  �R  S  ph  sO  r�%  �S  r"y  ��P  rfc ��P  rL �S   �O  �P  o�?  S  $S  ph  WL   s�B  NS  &�$  (  r\C  �NS  r?)  �SS   �J  �J  og6  fS  �S  ph  �M  x__s ^�  r^F  ^�+  vy�&  `uJ    ob  �S  �S  ph  LK   o�6  �S  �S  ph  �M  q__s �S  t^F  �+   �F  o�?  �S  T  ph  WL  r�%  �,   o);  T  3T  ph  3T  q__s 18T  t^F  1�+   �J  �F  o�<  KT  mT  ph  mT  q__s �rT  t^F  ��+   �J  �F  o{>  �T  �T  ph  �T  q__s ��T  t^F  ��+   �J  �F  o;  �T  �T  ph  3T  q__s �  t^F  �+   o�<  �T  U  ph  mT  q__s ��  t^F  ��+   oV>  U  AU  ph  �T  q__s y�  t^F  z�+   z�7   H^   �XU  �U  {h  �M  � |__s �]J  �|__n �H4  �}�N  -H   �~�N  9D 6H�2    �
7  �H�   ��U  �V  {h  �M  � ���  ��&  �H4  oD ��
 �
E  �D ��N  �H   �V  ~�N  �D �H�2   �6O  �H�  �>V  ~IO  E  I�B   �[O  �H	   �\V  ~iO  "E  �xO  �H
   �zV  ~�O  5E  �H4    ��M   X  I.   ��V  �V  ��M  � � �  �V  ��M  HE  �I   ~�M  gE �I   ��M  �I   ��M  �E     o�9  W  8W  ph  �M  tQ  �H4  vw�
 �
E  w8 �
E    �V7  0IN  �PW  pY  {h  �M  � |__i k�5  ��8�  ��&  m�5  �E ��
 n
E  �E �X�  �Nc z
E  F w �  {
E  �Y�  |�5  AF �wM  NIx�  {�W  ~�M  _F ~�M  �F  �WK  dI   X  ~eK  �F ~nK  G  �[M  jI   �6X  ~eM  G  ��M  �I   �UX  ~�M  +G  ��V  �I��  u�X  ~W  CG ~W  XG ���  �W  kG �*W  ��N  �I��  ��X  �O  �O  �O   } N  �I	   �~ON  �G ~CN  �G ~7N  �G ~.N  �G    �\N  FJ��  �RY  �jN  S���  �jN  S� N  vJ   ��ON  s� ��CN  P�7N  P�.N  S   �?M  OJ�  �~IM  �G     �A9  �J(  ��Y  �[  {h  �M  � |__s ~�  �|__n ~H4  ��(�  ��&  �H4  �G �8 �
E  H �6O  �JH�  �Z  ~IO  9H �K�B   ��O  �J	   �!Z  ~�O  WH  �`�  �[  �If ��B  jH �*W �H4  �H w_X ��B  ��R  �J   ��Z  ~�R  �H ~�R  �H  �x�  ��a ��B  �H ���  ��  I ��V  PK��  ��[  ~W  :I ~W  NI ���  �W  aI �*W  {I � N  YK��  �$[  ~ON  �I ~CN  �I ~7N  �I ~.N  �I  ��N  bK   �U[  ~O  �I ~O  �I ~O  �I  }�N  �K   �~O  
J ~O  /J ~O  NJ    Kr3    �HK�0    �07  �Kb  ��[  �`  {h  �M  � ���  ��&  Σ5  P��
 �
E  aJ ���  ��_ ��B  �J ��Z �qC  �J ���  �H4  {K �__r �1  CL �tN  �K �  ܏\  ~�N  �L ��N0   ~�N  ,M � N  �N�  �~ON  ?M ~CN  RM ~7N  eM ~.N  yM    �6O  �K@�  �\  ~IO  �M P�B   ��O  L	   ��\  ~�O  �M  �X�  �^  y�N ��F  ��P �H4  �M ��a �H4  �M �K_ ��B  <N �[O  L	   �7]  ~iO  eN  ���  n]  ���  
�  xN IOP�  pOi�  �O~�   ���  c^  ��d .]J  �\���  �]  �W_ &H4  �N M�3  P�B   �SN-   ^  ��P 6�
  �N }�O  dN   8��O  ~�O  �N ~�O  �N oN~�    ��O   N�  0~NP   O ~CP  FO ~8P  jO ~-P  �O ~"P  �O ~P  �O ~P  �O ~P   P   �xO  �O	   ��^  ~�O  P  �O��   ��V  CM0�  V1_  ~W  (P ~W  =P �0�  �W  PP �*W  ��N  PM`�  ��^  ~O  jP ~O  jP ~O  ~P  � N  iMx�  �~ON  �P ~CN  �P ~7N  �P ~.N  �P    ��V  �M��  M`  ~W  �P ~W  �P ���  �W  	Q �*W  � N  �M   ��_  ~ON  #Q ~CN  VQ ~7N  VQ ~.N  tQ  ��N  �M   ��_  ~O  �Q ~O  �Q ~O  �Q  } N  �N   ��ON  �CN  �7N  �.N     �[M  �M   O#`  ~eM  �Q  ��V  �M��  ��`  ~W  �Q ~W  �Q ���  �W  �Q �*W  ��N  �M   ��`  ~O  R ~O  R ~O  "R  } N  N	   �~ON  5R ~CN  5R ~7N  5R ~.N  HR    3M�3  �N�B  ;O�B  �O�B     �9   P�  �a  �d  {h  �M  � �__s &�  [R �__n &H4  S ���  ��&  )H4  �S ��
 @
E  ?T ��_ A�B  iT �tN  ]P��  3�a  ~�N  U �]P%   ~�N  GU � N  oP�  �~ON  [U ~CN  nU ~7N  �U ~.N  �U    �6O  �P0�  C�a  ~IO  �U �R�B   ��O  �P	   Cb  ~�O  �U  �H�  d  ��P G�B  �U �R'  TH4  �U ��V  /Qp�  q�b  ~W  *V ~W  ?V �p�  �W  SV �*W  � N  3Q��  ��b  ~ON  pV ~CN  pV ~7N  pV ~.N  �V  }�N  :Q   �~O  �V ~O  �V ~O  �V    ��O  R��  J'c  ~�O  �V ~�O  �V ~�O  �V R~�   ��V  0R��  id  ~W  W ~W  'W ���  �W  RW �*W  �W � N  >R��  ��c  ~ON  �W ~CN  �W ~7N  �W ~.N  �W  ��N  NR   ��c  ~O  
X ~O  
X ~O  X  }�N  �R
   �~O  2X ~O  WX ~O  vX    Q�3  �R�B   ��V  �Q �  9�d  ~W  �X ~W  �X � �  �W  �X �*W  � N  �Q�  ��d  ~ON  �X ~CN  �X ~7N  �X ~.N  �X  }�N  �Q   �~O  �X ~O  �X ~O  
Y    �WK  �R0�  /�d  ~eK  Y ~nK  <Y  �Q�0    �\N  �S  S+   �e  [e  �jN  � �
S!   ~jN  \Y � N  S   �~ON  pY ~CN  �Y ~7N  �Y ~.N  �Y    �tN  �\ 0S1   �we  �e  ��N  � �;S$   ~�N  �Y � N  CSP�  �~ON  �Y ~CN  �Y ~7N  Z ~.N  Z    o6   �e  �e  ph  �M   ��e  �[ pS  ��e  vf  ��e  � ��N  |Sp�  U+f  ~�N  *Z ��S �L  sT   UNf  �L  S��T ��S3TC  YT4C  �sT�T��   ��N  ��  �T
   ��f  �f  ~�N  �Z ��T�2   ��N  & �T7   ��f  �f  ��N  � ��T   ��N  S�TP�    z�6  �T`   ��f  g  {h  �M  � �Ti�  Ui�   ��7  @U8  �6g  Zi  {h  �M  � ��R ��  ����  �H4  ����  �W_ �H4  �Z ���  �H4  �Z �6O  RU��  ��g  ~IO  �Z xV�B   ��O  ZU	   ��g  ~�O  [  ���  ��P �H4  +[ ���  ��  u[ �9\ ��  �X��d �Zi  �\�__r �1  �[ �xO  mU	   �Ih  ~�O  �[  ��P  �U��  ��h  ~Q  �[ ~	Q  �\ ~�P  ] ~�P  B] ~�P  �] ~�P  (^ ~�P  H^ ��P   � V9   <i  ��N Zi  h^ ��a H4  �^ ��P  #V   2i  ~Q  �^ ~	Q  :_ ~�P  Y_ ~�P  l_ ~�P  �_ ~�P  �_ ~�P  �_ ~�P  �_  VVJ3   �UJ3  VJ3  sV�B     �9  �MR  5O �V[   �|i  j  �[R  � �dR  ���O  �V   1�i  ~�O  �_  ��V&   �dR  �~[R  ` ��V&   �qR  &` �R  �V�  :~<R  9` ~1R  ^` ~&R  s` �R  �~R  �`     �r9  �V`  �7j  �k  {h  �M  � � �  �a�  EqC  �` � X   zj  �Y�  H�9  �`  �6O  W@�  N�j  ~IO  �` @X�B   ��O  W	   N�j  ~�O  a  �X�  w�P T�B  ���  U�k  ��~�__r V1  a ���  WH4  Xa �p�  �k  �4 [�  ��~��R  <W��  \dk  ~�R  �a ~�R  �a ~�R  b ~�R  Hb ~�R  wb  ���  �W_ f�B  �b �WJ3    ��W!   �Y�  t�9  �b     iQ   �k  ��   zo8  @X�   ��k  m  {h  �M  ��Q  �5  ��@  �+  ���%  �4  ����  ��&  �5  � �tQ  WX   Fl  ��Q  ~�Q  �b  ���  m  �R �5  �b ��V  �X �  !�l  �W  ~W  c � �  �W  .c �*W  ��N  �X �  ��l  �O   �O   ~O  ]c  } N  �X	   ��ON  Q�CN  Q�7N  Q~.N  |c    �X�3   kXj    z�7  �X�  �)m  �p  {h  �M  � |__c ��5  ��8�  ��&  ��5  w �  �
E  �8 �
E  �c �X�  n  ��d ��F  �c �tN  �Xp�  ��m  ~�N  �c � Z0   ~�N  �c � N  	Z��  �~ON  �c ~CN  d ~7N  %d ~.N  9d    YMR  %Y�k   �wM  ;Y   �;n  ��M  �S�  ��M  �h�   �?M  IY   �Zn  ~IM  Ld  ��K  MY   ��n  ~�K  dd ~�K  wd  ��V  �Y��  �So  ~W  �d ~W  �d ���  �W  �d �*W  �d ��N  �Y   ��n  �O  �O  �O   � N  �Y��  �%o  ~ON  e ~CN  e ~7N  e ~.N  ?e  }�N  �Z   �~O  ]e ~O  �e ~O  �e    �?M  �Y   �ro  ~IM  �e  ��K  �Y   ��o  ~�K  �e ~�K  �e  ���  �o  �� ��4  �d�?M  �Y��  ��o  ~IM  �e  ��M  �Y   ��o  ~�M  f  �Zg   ��V  0Z`   ��p  ~W  3f ~W  Gf �0Z`   �W  Zf �*W  tf � N  9Z�  �{p  ~ON  �f ~CN  �f ~7N  �f ~.N  �f  ��N  BZ   ��p  ~O  �f ~O  �f ~O  �f  }�N  tZ   �~O  g ~O  (g ~O  Gg    fYg    �8  �Z  ��p  �r  {h  �M  ��Q  ��5  ��@  ��+  ���+  �� �  �8w  ��   Zg ��&  ��5  � ���  �
E  �g �[O  �Z   ��q  ~iO  �g  �tQ  [@�  ��q  ��Q  ��Q  �  ��N  ![X�  ��q  ~�N  �g K[�2   ���  ��b �qC  #h ��%  ��4  �S��N ��5  gh ���  5r  �R ��5  i �[�3   ��O  �[	   �Tr  ~�O  3i  �tN  �[+   ��r  ~�N  Fi ��[%   ~�N  pi � N  �[��  �~ON  �i ~CN  �i ~7N  �i ~.N  �i    E\�k  �\MR  �\MR     z>8  �\�   ��r  �s  {h  �M  ��%  �5  ���+  ����  ��&  	�5  � ��N  �\��  
Us  ~�N  �i ]�2   �tQ   ]   	{s  ��Q  ~�Q  �i  �tN  ]�  �s  ~�N  $j �`]'   ��N  S� N  i] �  ȆON  R�CN  P�7N  s4�.N  S   :]�k    ��8  �]�  �t  iv  {h  �M  � �ȱ  �iv  ��@�  �a�  �qC  Bj �Q �cJ  �j ��N  �]   �nt  ~�N  �j �]�2   �6O  �]`�  ��t  ~IO  Hk 9_�B   �[O  �]	   ��t  ~iO  [k  �6O  ^   ��t  ~IO  nk  ��O  ^	   ��t  ~�O  �k  ��O  3^	   �u  ~�O  �k  ��Q  Z^   �7u  ��Q  ~�Q  �k  ��^T   �u  �K_ ��B  �k �R  �^x�  ��u  ~<R  �k ~1R   l ~&R  5l ~R  Hl ~R  ul  /_��   ��V  �^&   �Lv  ~W  �l ~W  �l ��^&   �W  �l �*W  ��N  �^   �v  ~O  �l ~O  �l ~O  �l  } N  �^   �~ON  �l ~CN  �l ~7N  �l ~.N  m    �]C  �]4C  �^j    ZG  ��V  < @_u   ��v  }w  ~W  m ~W  6m ���  �W  Um �*W  �m � N  X_   ��v  ~ON  �m ~CN  Fn ~7N  Fn ~.N  n  ��N  �_   �!w  ~O  �n ~O  �n ~O  �n  ��N  �_   �Rw  ~O  �n ~O  �n ~O  �n  } N  �_   ��ON  �CN  �7N  �.N     z�:  �_   ��w  �w  {h  �w  �  �J  z�:  �_
   ��w  �w  �h  3T  o }�N  �_
   	~�N  %o ��_�2    z�:  �_
   �x  :x  �h  �w  =o }�N  �_
   ~�N  Qo ��_�2    zP<  �_   �Qx  ^x  {h  ^x  �  �J  zo<   `
   �zx  �x  �h  mT  io }�N   `
   �~�N  }o �
`�2    z�<  `
   ��x  �x  �h  ^x  �o }�N  `
   �~�N  �o �`�2    z�=   `   �y  y  {h  y  �  �J  z>  0`
   �7y  jy  �h  �T  �o }�N  0`
   e~�N  �o �:`�2    z7>  @`
   ��y  �y  �h  y  �o }�N  @`
   k~�N  p �J`�2    z�6  �`  ��y  �|  {h  �M  � ���  �|  ���  �qC  p ��N  �`   �z  ~�N  tp �`�2   ���  �|  	�_ �|{  
pe �iJ   ��_ Hz  dz  Mz  "z  Xz  e^z  "z   ��_ �uz  �z  ph  ~z  Mz  re �iJ   ��_ ��z  �z  ph  ~z  p#  �F   ��z  V P`K   ��z  ��z  � ��V  m`��  �q{  �W  �W  P���  �W  p,80.��*W  ��N  x`   �>{  �O   �O   �O  P } N  �`	   ��ON  R�CN  R�7N  R�.N  P   k`�f    ���  �"z  �\�dz  �`   ��{  ~�z  �p ~uz  >q  ��z  �`C   �}|  ~�z  mq ��V  �`�  �s|  ~W  �q ~W  �q ��  �W  �q �*W  ��N  �`   �<|  ~O  �q ~O  �q ~O  �q  } N  a	   �~ON  �q ~CN  �q ~7N  �q ~.N  �q    �`�f   �(�  �|  ��|  XaҲ  `a�2  ha�  �a�   �`j  qaҲ  ya�  ��a a�2   �a��     . �|  �  �|  e�|  o)6  }  %}  ph  �M  p#  �F   �}  kg �a6   �A}  {}  �}  � �L  �a@�  �k}  �L  ��a �a�y  ��a o�.  �}  �}  ph  �L  p#  �F  p�!  �}   �J  o
:  �}  �}  ph  3T  p#  �F  p�!  �}   �J  ��}  8d �a�   ��}  ~  ��}  � ��}  ��{}  �a`�  �8~  ~�}  r ~�}  Mr $b�?   ��L  hb   �`~  ��L  v���L  S �9bIb�?  �bbb��   ��}  hb �b�   ��~  D  ��}  � �S  �bI   ��~  ~S  �r ��b �{}  �b   ��~  ��}  ,	�~�}  �r �b�?   �6L  5c   �%  �DL  s� ��Ec �cc�?  �/cMc��   o�;  R  n  ph  mT  p#  �F  p�!  n   �J  �D  �T Pc�   ��  �  �R  � �d  ��bL  _cx�  t�  ~�L  s ~pL  Gs yc�?   �M  �c   t�  �0M  v��M  S ��c�c�?  ��c�c��   �D  S �c�   �5�  ׀  �R  � �S  �cI   tc�  ~S  }s ��c �bL  5d   t��  ��L  ~pL  �s Ld�?   �6L  �d   t��  �DL  s� ���d �ddmd�?  ��d�d��   �>  o�>  �  �  ph  �  p#  �F  p�!  �   ׀  �J  o\=  �  ;�  ph  �T  p#  �F  p�!  ;�   �J  ��  �d �d�   �\�  I�  ��  � �1�  ��݀  �d��  '�  ~��  �s ~�  \t �{}  �d"   	?Ɓ  ~�}  �t ~�}  \t �d�?   �bL  �d   	?��  ~�L  �t ~pL  Pu �d�?   }�L  Ue   	?~�L  �u ~�L  �u   �/e?e�?  le��  �ue��e�e��   ��  �b �e  �e�  a�  ��  � �S  �eI   '��  ~S  �u ��e �݀  �e6   '�  ~��  v ~�  Fv �{}  �e    	?�  ��}  ~�}  Fv f�?   }bL  f   	?~�L  |v ~pL  �v f�?    �6L  zf   '<�  �DL  s� ���f �:fCf�?  �df�wf�f��   �XS  �^ �f�   �}�  �  �fS  � �oS  ��zS  ���f7   �  ��S  �v ��N  �f   a׃  ~�N  w �f�2   ��N  �f   d��  ~�N  Rw �f�2   �f;2   ���  ~oS  |w ~zS  �w ~fS  �w ���  ��S  ��V  �f��  lل  ~W  �w ~W  �w ���  �W  #x �*W  ��N  g��  ���  ~O  _x ~O  _x ~O  sx  } N  g	   �~ON  �x ~CN  �x ~7N  �x ~.N  �w    �f�N  ^g�y     ��S  �O �g   �
�  C�  ��S  � ~�S  �x ��S  ���gXS  �� � ���  �T  �P �g\   �_�  \�  �T  � �T  ��&T  ���Q  �g�  3��  ��Q  ~�Q  �x  ��S  �g �  3څ  ~�S  �x ~�S  !y ~�S  Ay �gXS   �8�  Q�  ~T  �y �&T  �~T  �y ��S  �gP�  4��S  ~�S  �y ��M  �gh�  �E�  �N  ~	N  �y  ��g@    ��g@   �=T  Z �g\   �x�  u�  �KT  � �TT  ��`T  ���Q  �g��  ���  ��Q  ~�Q  z  ��S  �g��  ��  ~�S  +z ~�S  Rz ~�S  rz hXS   ���  j�  ~TT  �z �`T  �~KT  �z ��S  5h��  ���S  ~�S  �z ��M  5h��  �^�  �N  ~	N  {  �Lh@    �0h@   �wT  �W Ph\   ���  h�  ��T  � ��T  ���T  ���S  Xh��  ��  ��S  �~�S  ={ ~�S  ]{ khXS   ��  ]�  ~�T  �{ ��T  �~�T  �{ ��S  �h(�  ���S  ~�S  �{ ��M  �h@�  �Q�  �N  ~	N  	|  ��h@    ��h@   ��T  �` �h\   ���  P�  ��T  � ��T  ���T  ���Q  �hX�  ň  ��Q  ~�Q  (|  �p�  <�  ~�T  G| ��T  �~�T  [| ��S  �h��   ��S  ~�S  z| ��M  �h��  �0�  �N  ~	N  �|  �i@    �hXS  ��h@   ��T  4P i\   �l�  8�  ��T  � ��T  ��U  ���Q  i��  ���  ��Q  ~�Q  �|  ���  $�  ~�T  �| �U  �~�T  �| ��S  Ui��  ���S  ~�S  
} ��M  Ui �  ��  �N  ~	N  )}  �li@    -iXS  �Ni@   �U  �U pi\   �T�  ��  �U  � �(U  ��4U  ���  �  ~(U  H} �4U  �~U  \} ��S  �i0�  }��S  ~�S  {} ��M  �iH�  �ڊ  �N  ~	N  �}  ��i@    �iXS  ��i@   o�>  �  0�  ph  �  p#  �F  p�!  0�  t(  	4QK   �J  �.  o�.  I�  p�  ph  �L  p#  �F  p�!  p�  r(  	]5�   �J  o}=  ��  ��  ph  �T  p#  �F  p�!  ��  q__s 3�  t^F  4�+   �J  �u�  `] �i7  �؋  ��  ���  � ���  ����  ����  ����  �i`�  5��  �#�   ~�  �} ~�  3~ �;�  �i"   	5b�  �d�   ~[�  �~ ~I�  3~ j�?   ��L  j   	5��  ��L   ~�L   ~�L  � j�?   }�L  �j   	5~�L  � ~�L  �   �U  bj��  8�  ~4U  � ~(U  S� ~U  �� ��j   l�  ~(U  ـ ~4U  �� ~U  � ��S  �j��  }~�S  D� ~�S  X� ��M  �j   �a�  ~N  D� ~	N  k�  �j@    njXS  �j@   �Oj_j�?  �j��  ��j��jk��   o�=  ��  �  ph  �T  p#  �F  p�!  �  q__s B�  t^F  C�+   �J  �F  ���  �X k7  ��  �  ���  � �͍  ��֍  ���  ����  k��  D��  �#�   ~�  � ~�  �� �;�  k"   	5��  �d�   ~[�  R� ~I�  �� Ak�?   ��L  Ak   	5׎  ��L   ~�L  ΂ ~�L  J� ]k�?   }�L  l   	5~�L  �� ~�L  ΃   �wT  �k��  G�  ~�T  � ~�T  � ~�T  Q� ��S  �k��  �e�  ~�S  � ~�S  � ~�S  �� �kXS   ��k   �  ~�T  �� ~�T  � ~�T  =� ��S  �k�  �~�S  h� ~�S  |� ��M  �k   �؏  ~N  h� ~	N  ��  �k@    �k@   ��k�k�?  $l��  �-l�?lGl��   �u�  �c PlV  �7�  �  ���  � ���  ����  ��S  \lI   5w�  ~S  �� �el ���  �l6   5�  �#�   ~�  � ~�  Z� �;�  �l    	5ڐ  �d�   �[�  ~I�  Z� �l�?   }�L  �l   	5~�L  �� ~�L  ӆ ~�L  �� �l�?    �U  m �  8ё  ~4U  j� ~(U  �� ~U  ڇ �@m   ��  ~(U  (� ~4U  H� ~U  h� ��S  Bm8�  }~�S  �� ~�S  �� ��M  Jm   ���  ~N  �� ~	N  ��  Wm@    mXS  +m@   �6L  �m   5��  �DL  s� ���m ��lm�?  �xm��m�m��   ���  o^ �mV  �9�  P�  ���  � �֍  ���  ��S  �mI   Dy�  ~S  Έ ��m ���  n6   D�  �#�   ~�  E� ~�  �� �;�  n    	5ܒ  �d�   �[�  ~I�  �� #n�?   }�L  %n   	5~�L  މ ~�L  �� ~�L  &� ;n�?    �wT  cnP�  G�  ~�T  �� ~�T  ͊ ~�T  � ��S  cnp�  �|�  ~�S  �� ~�S  ͊ ~�S  S� tnXS   ��n   ��  ~�T  �� ~�T  ы ~�T  � ��S  �n��  �~�S  � ~�S  0� ��M  �n   ��  ~N  � ~	N  C�  �n@    �n@   �6L  �n   D+�  �DL  s� ���n �Zncn�?  ��n��no��   o�;  ^�  ��  ph  mT  p#  �F  p�!  ��  q__s ��  t^F  ��+   �J  �P�  �O o�   ���  8�  �^�  � �p�  ��y�  ����  ��bL  o��  ��  ~�L  W� ~pL  ƌ 9o�?   ��T  ^o��  ��  ~U  � ~�T  W� ~�T  �� ��Q  ^o��  �`�  ~�Q  ݍ ~�Q  �  ��o   ޕ  ~�T  � ~U  � ~�T  1� ��S  �o��  �~�S  \� ~�S  p� ��M  �o   �ӕ  ~N  \� ~	N  ��  �o@    qoXS  �o@   �M  �o   ��  �0M  v��M  S �No^o�?  ��o�o��   o�;  F�  z�  ph  mT  p#  �F  p�!  z�  q__s ��  t^F  ��+   �J  �F  �8�  �f �o�   ���  V�  �F�  � �X�  ��a�  ��m�  ��bL  �o�  ���  ~�L  �� ~pL  � p�?   �=T  >p �  ��  ~`T  _� ~TT  �� ~KT  Ϗ ��Q  >p@�  �M�  ~�Q  � ~�Q  _�  ��S  Gp   ���  ~�S  1� ~�S  �� ~�S  y� SpXS   ��p   �  ~TT  א ~`T  �� ~KT  � ��S  �pX�  �~�S  B� ~�S  V� ��M  �p   ���  ~N  B� ~	N  i�  �p@    lp@   �M  �p   �7�  �0M  v��M  S �.p>p�?  ��p�p��   o+:  d�  ��  ph  3T  p#  �F  p�!  ��  q__s ��  t^F  ��+   �J  �V�  �e �p�   ���  >�  �d�  � �v�  ���  ����  ��{}  �pp�  ��  ~�}  }� ~�}  � q�?   ��T  )q��  ���  ~�T  E� ~�T  }� ~�T  �� ��Q  )q��  f�  ~�Q  � ~�Q  E�  �`q   �  ~�T  � ~�T  7� ~�T  W� ��S  bq��   ~�S  �� ~�S  �� ��M  jq   �ٙ  ~N  �� ~	N  ��  wq@    <qXS  Uq@   ��L  �q   ��  ��L  v���L  S �q)q�?  ��q�q��   oV:  L�  ��  ph  3T  p#  �F  p�!  ��  q__s ���  t^F  ��+   �J  �F  �>�  Ma �q�   ���  \�  �L�  � �^�  ��g�  ��s�  ��{}  �q��  ���  ~�}  �� ~�}  ,� �q�?   �T  	r��  ��  ~&T  �� ~T  �� ~T  �� ��Q  	r�  3S�  ~�Q  C� ~�Q  ��  ��S  r   3��  ~�S  W� ~�S  �� ~�S  �� rXS   �Pr   �  ~T  �� ~&T  � ~T  =� ��S  Rr(�  4~�S  h� ~�S  |� ��M  Zr   � �  ~N  h� ~	N  ��  gr@    7r@   ��L  �r   �=�  ��L  v���L  S ��q	r�?  ��r�r��   �P�  �` �r   �x�  �  �^�  � �y�  ����  ��S  �rI   ���  ~S  �� ��r �bL  �r   ��  ��L  ~pL  � s�?   ��T  -s@�  �ϝ  ~U  s� ~�T  �� ~�T  � ��Q  -s`�  �>�  ~�Q  1� ~�Q  s�  �ps   ��  ~�T  E� ~U  e� ~�T  �� ��S  rsx�  �~�S  �� ~�S  Ę ��M  zs   ���  ~N  �� ~	N  ט  �s@    @sXS  Ys@   �6L  �s   ���  �DL  s� ���s �$s-s�?  ��s�s��   �8�  T �s   �1�  ��  �F�  � �a�  ��m�  ��S  �sI   �q�  ~S  � ��s �bL  t   ���  ��L  ~pL  b� ,t�?   �=T  Mt��  ���  ~`T  �� ~TT  � ~KT  +� ��Q  Mt��  ���  ~�Q  y� ~�Q  ��  ��S  Vt   �1�  ~�S  �� ~�S  � ~�S  ՚ btXS   ��t   ��  ~TT  3� ~`T  S� ~KT  s� ��S  �t��  �~�S  �� ~�S  �� ��M  �t   ���  ~N  �� ~	N  ś  �t@    {t@   �6L  �t   ���  �DL  s� ���t �DtMt�?  ��t�t��   �V�  g �t   ��  ��  �d�  � ��  ����  ��S  �tI   �[�  ~S  ٛ ��t �{}  5u   ���  ��}  ,	�~�}  P� Su�?   ��T  tu��  �y�  ~�T  �� ~�T  � ~�T  � ��Q  tu �  �  ~�Q  g� ~�Q  ��  ��u   f�  ~�T  {� ~�T  �� ~�T  �� ��S  �u�   ~�S  � ~�S  �� ��M  �u   �[�  ~N  � ~	N  �  �u@    �uXS  �u@   �6L  �u   ���  �DL  s� ���u �kutu�?  ��u v��   �>�  �N  v   �ۡ  ��  �L�  � �g�  ��s�  ��S  vI   ��  ~S  !� �v �{}  Uv   �P�  ��}  ,	�~�}  �� sv�?   �T  �v0�  �j�  ~&T  � ~T  )� ~T  a� ��Q  �vP�  3��  ~�Q  �� ~�Q  �  ��S  �v   3�  ~�S  ß ~�S  )� ~�S  � �vXS   ��v   `�  ~T  i� ~&T  �� ~T  �� ��S  �vh�  4~�S  Ԡ ~�S  � ��M  �v   �U�  ~N  Ԡ ~	N  ��  �v@    �v@   �6L  w   ���  �DL  s� ��w ��v�v�?  �w w��   zN;   w=   �ǣ  1�  {h  3T  � ��S  Bw��  F'�  ��S  ~�S  � ��M  Hw   ��  �N  ~	N  "�  Uw@   1w�y   z�<  `w=   �H�  ��  {h  mT  � ��S  �w��  ���  ��S  ~�S  6� ��M  �w   ���  �N  ~	N  I�  �w@   qw�y   z�>  �w=   �ɤ  3�  {h  �T  � ��S  �w��  �)�  ��S  ~�S  ]� ��M  �w   ��  �N  ~	N  p�  �w@   �w�y   �}  �N �w=   �O�  ��  �}  � �}  �w(   ܩ�  ~}  �� �L  �w   ܙ�  ~L  �� �x �w�y  ��w �x�   o*<  ¥  ޥ  ph  mT  p#  �F  p�!  ޥ   �J  ���  I`  x[   ���  ��  �¥  � �ԥ  ��}  =x*   �c�  ~}  ¡ �L  Ux   �S�  ~L  �� �gx Jx�y  �Ux }M  gx   �~0M  $� ~M  I�   o�:  ��  ��  ph  3T  p#  �F  p�!  ��   �J  ���  �W �x[   �Ҧ  Z�  ���  � ���  ��}  �x*   �6�  ~}  h� �L  �x   �&�  ~L  �� ��x �x�y  ��x }�L  �x   �~�L  ʢ ~�L  �   ���  @^ �xX   �v�  �  �¥  � �}  �x��  �ѧ  ~}  � �L  y��  ���  ~L  ]� �%y y�y  �y �6L  y��  ��DL  �8y  ���  cU PyX   ��  ��  ���  � �}  hy�  �g�  ~}  �� �L  �y0�  �W�  ~L  � ��y uy�y  ��y �6L  �yH�  ��DL  ��y  o?  ��  ��  ph  �  p#  �F  p�!  ��   �J  o�=  è  ߨ  ph  �T  p#  �F  p�!  ߨ   �J  ���  �d �y�   � �  ө  �è  � �ը  ��}  �yh�  Rd�  ~}  4� �L  �y   �T�  ~L  q� �z �y�y  ��y }��  z2   R~��  �� ~��  �� �M  !z   	;��  ~0M  ڤ ~M  ��  }�L  1z   	;~�L  $� ~�L  I�    ���  n\ Pza   ��  ��  �¥  � ���  XzL   ���  ~¥  h� �}  hz*   �h�  ~}  �� �L  �z   �X�  ~L  �� ��z uz�y  ��z }6L  �z   �~DL  ܥ ��z  ��z�   ���  nS �za   ���  U�  ���  � ���  �zL   �J�  ~��  � �}  �z*   �)�  ~}  :� �L   {   ��  ~L  j� �{ �z�y  � { }6L  {   �~DL  �� �${  �1{�   ���  hV P{_   �q�  �  �è  � �}  o{��  R̫  ~}  Φ �L  �{��  ܼ�  ~L  � ��{ |{�y  ��{ �6L  �{��  R�DL  ��{  ���  \ �{h   ��  ��  �è  � ���  �{S   R��  ~è  a� �}  �{*   R��  ~}  �� �L  |   �p�  ~L  �� �| �{�y  �| }6L  |   R~DL  է �+|  �8|�   �U  =��   �  ��   >��  �B  ?��  ��  E�   �  �B   F�  �C  G�  �e  H�  �8  I�  ��  J�  �

  X8�   �  ��  Y8�  ��
  Z8�  ��   `d�  �  ��  fv�   �  ��  gv�  ��  hv�  ��  n��   �  ��	  o��  ��  p��  �H  vέ   	  �`  wέ  �w  xέ  �   yέ  �~  �     �   ��  ��  ��  �  ��  ��   ��  ��  ��  ��	  ��  ��  �g�     �  �g�  �  �g�  ��  �g�  ��  ���   *  ��  ���  ��  ���  ��  ���  �m  �ٮ   5  �	  �ٮ  �2	  �ٮ  ��  �ٮ  �9  �ٮ  �[  ��   @  �J  ��  ��  ��  �7  ��  ��  �X�   K  �I	  �X�  �$	  �X�  ��   ���   V  �N  ���  �p  ���   a  ��  ���  �:  ���  ��  £�  �d   ã�  ��  ��   l  �  ��  ��  ��  ��	  ��   w  ��  ��  �  �4�   �  ��  �4�  ��  �4�  ��  �4�  �+  �m�   �  ��  �m�  ��   �m�  �  陰   �  ��
  ꙰  ��  뙰  �  �Ű   �  �   �Ű  �F  �Ű  ��  ��   �  ��  ��  ��  ��  �D  O�   �  ��  P�  �1  Q�  ��  WI�   �  �^  XI�  ��  3h�   �  ��  4h�  ��   8��   �  ��  9��  �l	  =��  �  �N  >��  �^  ?��  �L  @��  �a  D߱  �  �B  E߱  ��	  F߱  �  G߱  �  H߱  �y  I߱  ��   2�   
  ��  !2�  ��B  �0  c�  /��  �  i�  �
   !�e  /�Ӫ  ~�  �   ��d  �  ��  �  �  �   ��O �O �  ��  �  �  7    �>  Y  Ҳ  �   ��  �  �  �   ��  ��  ��  /�1  �    �   y�  �p p �b �     �6 std " 1+  ++ 	S�S 
L��  Y�$ _[   @     ��  cn   H     �  g�   [     %  0@�5  �=  �W  �b  � 3  Fe  ��2  	�3  �=  �   
�5  
�5   �   eq �<-  �2  �   
�5  
�5   lt ��1  �2  
  
�5  
�5   ��  eF  �2  .  
�5  
�5  
W   �K  �9  W  H  
�5   �(  
!  �5  l  
�5  
W  
�5   1  �A  �5  �  
�5  
�5  
W   �5  �'  �5  �  
�5  
�5  
W   �3  �A  �5  �  
�5  
W  
�    +  :  �   �  
�5   �   �C   �P  �     
�5   �B  $6  �2  0  
�5  
�5   eof (�:  �   ?  ,N0  �   
�5    _� ��2  023  1H3  2^3  3t3  5�3  6�3  74  84  :3  ;�3  <�3  =�3  ?E4  @/4  B'3  C=3  DS3  Ei3  G�3  H�3  I4  J$4  L�3  M�3  N�3  O�3  QP4  R:4  v  6�  x  K�  �  MZ5   x  OX  c  �5  
Z5   �  Qw  v  |  �5   �  R  �  �  �5     T8  Z5  �  �   6   x  Z�  �  �5   x  \�  �  �5  
6   x  _�  �  �5  
�   x  c    �5  
6   �  p�  6  1  <  �5  
6   �  t�  6  T  _  �5  
6   �  {o  z  �5  �2   n	 ~%  �  �  �5  
6   �  ��  �2  �  �   6   �  �h  6  �   6    1   :1  �  �3  � �  �?  ��2  K  \�  Q+   �e  _W  ��  `�  �4  c6  �J  d$6  ��  qR  X  <6   ��  sh  s  <6  
B6   W  y�  �  <6  �2   �k h�< i�   �h  3    �  5O6  6|7  7�7  �J  pG!  !�B  @  �   "%  M5   #�B      �7  
M5  
B6   $�B     +  �7  �2   %�B  4  �7  
@    �e  y  &[V  Y  @  "�G  !�   <  x�  ��  z  �4  {*  �J  |6  �J  �,  `S  ��.  ~J  �G!  �J  �z#  �%  ��  �K  �@   I  �@  :!  ��7   %H  ��  �   '�3  2Y  '�G  7�5  't3  B�7  	x ��  (�'  ��O  �7  V  ��N  �2  `  f  �7   3  �o+  �2  }  �  �7   �P  ��O  �  �  �7   �M  ��P  �  �  �7   �,  �-  �  �  �7  
@   �+  ��R  M5  �  �  �7   3  �   M5      �7  
B6  
B6   �/  !�B  �7  ;  
@  
@  
B6   �O  �|6  N  Y  �7  
B6   )(  ��6  m  x  �7  
B6   *�   �-  M5  �  �  �7   +�1  o�*  M5  �  �7  
B6  
@    *�A  $n%  M5  �  �  �7   *�A  (�I  M5  �  �  �7  
M5   *"A  ,�%  �7  	  	  �7   *�1  2E)  �  2	  8	  �7   *�/  6;&  �  P	  V	  �7   )�>  :�>  j	  p	  �7   *S  A:2  @  �	  �	  �7  
@  
�5   )�#  K�(  �	  �	  �7  
@  
@  
�5   *9  S>$  @  �	  �	  �7  
@  
@   *-U  [�7  �2  
  
  �7  
�5   ,�5  d�-  ,
  
M5  
�5  
@   ,	1  m�P  L
  
M5  
�5  
@   ,�3  v\-  l
  
M5  
@  
 3   ,nU  ��-  �
  
M5  
�  
�   ,nU  �nG  �
  
M5  
�  
�   ,nU  ��   �
  
M5  
M5  
M5   ,nU  �IP  �
  
M5  
�5  
�5   �J  �rR  �2    
@  
@   )�=  ��H    4  �7  
@  
@  
@   )V  �)  H  N  �7   -�'  �D*  �7  .�0  �o  u  �7   /�0  ��  �  �7  
B6   .�0  ��  �  �7  
�7   .�0  ��  �  �7  
�7  
@  
@   .�0  ��  �  �7  
�7  
@  
@  
B6   .�0  �  $  �7  
�5  
@  
B6   .�0  �5  E  �7  
�5  
B6   .�0  �V  k  �7  
@  
 3  
B6   .�0   |  �  �7  
�7   .�0  �  �  �7  
�%  
B6   .�0  "�  �  �7  �2   0�  *,Q  �7  �  �  �7  
�7   0�  2�G  �7      �7  
�5   0�  =�%  �7  %  0  �7  
 3   0�  Mo_ �7  I  T  �7  
�7   0�  Y.c �7  m  x  �7  
�%   0S� f�&  �  �  �  �7   0S� q�>  �  �  �  �7   1end y<  �  �  �  �7   1end �6;  �  �  �  �7   0I ��$  �      �7   0I ��7  �  ,  2  �7   0��  �lC  �  K  Q  �7   0��  �CM  �  j  p  �7   0)^ �^\ �  �  �  �7   0%] ��a �  �  �  �7   0hf �*] �  �  �  �7   0wY �Je �  �  �  �7   0r ��R  @      �7   0�K  �r5  @  $  *  �7   0�3  �j=  @  C  I  �7   2�� ��  ^  n  �7  
@  
 3   2�� ��F  �  �  �7  
@   2be  VT �  �  �7   0I  v  @  �  �  �7   2�E  &|U  �  �  �7  
@   2�1  -�  �    �7   0�� 5�?  �2    "  �7   0�:  D�6  �  ;  F  �7  
@   0�:  UW  �  _  j  �7  
@   1at k
/  �  �  �  �7  
@   1at ��7  �  �  �  �7  
@   0��  ��O �  �  �  �7   0��  �}Y �  �  �  �7   0�G  �@\ �      �7   0�G  �e �  &  ,  �7   0�F  ��/  �7  E  P  �7  
�7   0�F  �k:  �7  i  t  �7  
�5   0�F  ��H  �7  �  �  �7  
 3   0�F  �x` �7  �  �  �7  
�%   0@  �A:  �7  �  �  �7  
�7   0@  ��1  �7  �    �7  
�7  
@  
@   0@  ��D  �7  '  7  �7  
�5  
@   0@  ��*  �7  P  [  �7  
�5   0@  �6  �7  t  �  �7  
@  
 3   0@  �] �7  �  �  �7  
�%   2�G  -aN  �  �  �7  
 3   0�3  <b*  �7  �  �  �7  
�7   0�3  Ipf �7      �7  
�7   0�3  ^ 2  �7  )  >  �7  
�7  
@  
@   0�3  n�=  �7  W  g  �7  
�5  
@   0�3  z�T  �7  �  �  �7  
�5   0�3  � @  �7  �  �  �7  
@  
 3   0�3  ��a �7  �  �  �7  
�%   2� ��E  �    �7  
�  
@  
 3   2� ��V   '  �7  
�  
�%   0� �\+  �7  @  P  �7  
@  
�7   0� �u>  �7  i  �  �7  
@  
�7  
@  
@   0� |=  �7  �  �  �7  
@  
�5  
@   0� "�@  �7  �  �  �7  
@  
�5   0� 9k<  �7  �    �7  
@  
@  
 3   0� K�'  �  !  1  �7  
�  
 3   0bL  d�R  �7  J  Z  �7  
@  
@   0bL  t�2  �  s  ~  �7  
�   0bL  �L&  �  �  �  �7  
�  
�   2H�  �M\ �  �  �7   0�%  �9F  �7  �  �  �7  
@  
@  
�7   0�%  �|<  �7  	  (  �7  
@  
@  
�7  
@  
@   0�%  ��T  �7  A  [  �7  
@  
@  
�5  
@   0�%  ��A  �7  t  �  �7  
@  
@  
�5   0�%  b>  �7  �  �  �7  
@  
@  
@  
 3   0�%  3%  �7  �  �  �7  
�  
�  
�7   0�%  'V7  �7      �7  
�  
�  
�5  
@   0�%  <�+  �7  6  K  �7  
�  
�  
�5   0�%  Q'S  �7  d  ~  �7  
�  
�  
@  
 3   0�%  vj.  �7  �  �  �7  
�  
�  
M5  
M5   0�%  ��9  �7  �  �  �7  
�  
�  
�5  
�5   0�%  �C  �7  �    �7  
�  
�  
�  
�   0�%  �>/  �7  0  J  �7  
�  
�  
�  
�   0�%  �b �7  c  x  �7  
�  
�  
�%   *�?  ��&  �7  �  �  �7  
@  
@  
@  
 3   *�1  �O  �7  �  �  �7  
@  
@  
�5  
@   ,)  �z-  M5     
@  
 3  
B6   +E  �3J  M5  $  
@  
 3  
B6   0�5  �)  @  =  R  �7  
M5  
@  
@   2n	 @D  g  r  �7  
�7   0W�  �6  �5  �  �  �7   0�A  %�A  �5  �  �  �7   0��  ,Z5  k  �  �  �7   0�(  <;  @  �  �  �7  
�5  
@  
@   0�(  I�%  @    &  �7  
�7  
@   0�(  X�5  @  ?  O  �7  
�5  
@   0�(  i^   @  h  x  �7  
 3  
@   0�(  v�S  @  �  �  �7  
�7  
@   0�(  �K  @  �  �  �7  
�5  
@  
@   0�(  �o?  @  �  �  �7  
�5  
@   0�(  �J5  @    !  �7  
 3  
@   0NW  ��Q  @  :  J  �7  
�7  
@   0NW  ��I  @  c  x  �7  
�5  
@  
@   0NW  ��,  @  �  �  �7  
�5  
@   0NW  ��;  @  �  �  �7  
 3  
@   0�S  ��I  @  �  �  �7  
�7  
@   0�S  T?  @    !  �7  
�5  
@  
@   0�S  05  @  :  J  �7  
�5  
@   0�S  $S:  @  c  s  �7  
 3  
@   0�>  2hL  @  �  �  �7  
�7  
@   0�>  CUB  @  �  �  �7  
�5  
@  
@   0�>  Q�2  @  �  �  �7  
�5  
@   0�>  b�K  @      �7  
 3  
@   0�4  qT  @  5  E  �7  
�7  
@   0�4  ��K  @  ^  s  �7  
�5  
@  
@   0�4  ��5  @  �  �  �7  
�5  
@   0�4  �N.  @  �  �  �7  
 3  
@   0U+  �)  �  �  �  �7  
@  
@   0��  �!1  �2      �7  
�7   0��  ��T  �2  +  @  �7  
@  
@  
�7   0��  ��O  �2  Y  x  �7  
@  
@  
�7  
@  
@   0��  	;.  �2  �  �  �7  
�5   0��  (	�B  �2  �  �  �7  
@  
@  
�5   0��  C	�,  �2  �  �  �7  
@  
@  
�5  
@   �  w  �  3�q �M5  :   �  �,  
�,  
�,  
B6  
0    3�q �M5  c   �  �,  
�,  
�,  
B6   4�) {M5  �   ß  M5  
M5  
M5  
B6  
H    3E) �M5  �   �  M5  
M5  
M5  
B6  
0    3�) �M5  �   �  M5  
M5  
M5  
B6   4<�  {M5      ß  �5  
�5  
�5  
B6  
H    3��  �M5  B    �  �5  
�5  
�5  
B6  
0    3<�  �M5  k    �  �5  
�5  
�5  
B6   k  5�q {�n M5  �    ß  �,  
�,  
�,  
B6  
H    {* ��   �    f�  M5  �7  
M5  
M5  
B6   �  ��   �    f�  �5  �7  
�5  
�5  
B6   /t �!  +!   f�  �,  �7  
�,  
�,  
B6    !T   3  6�E  �   6�F  �   �&  az#  a(   7I�  i�.   �s n�.  ��  o6(  � pA(  �4  qL(  �J  y�!  �!  \8   8�J  �!  �!  \8  
g!   �J  ��!  �!  \8  
b8   WC  �v g!  �!  "  h8   *  ��u �!  "  "  h8   Ư  �ah !  7"  ="  h8   �F  �|n n8  U"  ["  \8   �F  ��m G!  s"  ~"  \8  
�2   a�  �6s n8  �"  �"  \8   a�  ��r G!  �"  �"  \8  
�2   (*  �l G!  �"  �"  h8  
s!   �F  �Pw n8  �"  #  \8  
s!   �O  ��t G!  #  (#  h8  
s!   0 I  �i n8  A#  L#  \8  
s!   0�:  �h �!  e#  p#  h8  
s!    {�  �.   �7  a�%  �'   7I�  i�,   �s n�,  ��  o�'  � p�'  �4  q�'  �J  y�#  �#  D8   8�J  �#  �#  D8  
�#   �J  �$  $  D8  
J8   WC  ��s �#  .$  4$  P8   *  �#r �#  L$  R$  P8   Ư  �n �#  j$  p$  P8   �F  �gx V8  �$  �$  D8   �F  �$x z#  �$  �$  D8  
�2   a�  �bl V8  �$  �$  D8   a�  �l z#  �$  �$  D8  
�2   (*  �^v z#  
%  %  P8  
�#   �F  �p V8  -%  8%  D8  
�#   �O  �Ai z#  P%  [%  P8  
�#   0 I  �v V8  t%  %  D8  
�#   0�:  rr �#  �%  �%  P8  
�#    {�  �,   �  Qf /�&  �J  6�5  t :�%   �e  5W  �x ;�%  `S  7�5  9�w >	&  &  88  
�%  
�%   �w B)&  /&  88   r G�i �%  G&  M&  >8   S� K�m �%  e&  k&  >8   :end O;u �%  �&  �&  >8   ;_E  3   <S +�  ד  ��&  �q  �n   ��  ��  � �M5  �4  �6   {�  M5   �u v'   |t �5   �t �5   �m �2   !np kJ'  �&   *V�  nzu �2  0'  @'  8  
8  
8   ;_Tp �5   '  �k  ��'  �q  �n   ��  ��  � ��5  �4  �$6   {�  �5   �%  qk ��'  �q  ��,  ��  ��,  � ��,  �4  ��,   {�  �,   �o v%(  $�J  �'  �'  ~=    �#  n   ;_Tp  3   �.  �2   �?  M5   �   6   z#  �g �a(  ��  ��.  � �/  �4  ��.   {�  �.   �w v�(  $�J  z(  �(  �=    �#  n   ;_Tp  3   �.  �2   �?  �5   �   $6   G!  4}�  ��2  �(  ;_Tp  3  
B6  
B6   4ͳ  �H>  �(  ;_Tp �2  
H>  
H>   46o ɢ'  )   8�  �,  
@B   4�j Z�'  ?)   ��  �,  
�,  
�,  
n    4�j r�'  b)   f�  �,  
�,  
�,   4P* ɧ&  �)   8�  M5  
�7   4�% Z�&  �)   ��  M5  
M5  
M5  
n    4�% r�&  �)   f�  M5  
M5  
M5   4�  �['  �)   8�  �5  
8   4z�  Zf'  *   ��  �5  
�5  
�5  
n    4|�  rf'  4*   f�  �5  
�5  
�5   �h �j �  n*   !T   3   �E  �    �F  �  
�5  
�7   �h ��o �  �*   !T   3   �E  �    �F  �  
 3  
�7   �h P	Um �  �*   !T   3   �E  �    �F  �  
�7  
�7   =	[ 
O�*   8   	��  N)�  
+  
�5  > 	� H� +  
�5   ?�p ?]u 
�5    $   	E�2  �  $,W  -�  K  :�,  �e  =W  � ?M5  "  @�5  �4  A6  �J  B$6  �A  O�+  �+  *6   �A  Q�+  �+  *6  
06   �A  V�+  �+  *6  �2   �
 Y51  i+  �+  ,  66  
�+   �
 ]�R  u+   ,  +,  66  
�+   � c?  i+  C,  S,  *6  
]+  
�5   _ m.   g,  w,  *6  
i+  
]+   �3  q89  ]+  �,  �,  66   ;_Tp  3   Q+  @ZD  ��.  AF�  �M5   B�q  ��&  B��  ��&  B�4  ��&  B� ��&  .��  �-  
-  �7   /��  �-  &-  �7  
�7   0*  ��}  �,  ?-  E-  	8   0Ư  �?s  �,  ^-  d-  	8   0�F  �Ϭ  8  }-  �-  �7   0�F  ��  �,  �-  �-  �7  
�2   0a�  �
�  8  �-  �-  �7   0a�   ��  �,  �-  �-  �7  
�2   0�:  ,�  �,  .  .  	8  
�,   0�F  		n  8  '.  2.  �7  
�,   0(*  ��  �,  K.  V.  	8  
�,   0 I  h�  8  o.  z.  �7  
�,   0�O  7k  �,  �.  �.  	8  
�,   0WC  ]�  �7  �.  �.  	8    {�  M5   �  �   @8E  ��0  AF�  ��5   B��  �f'  B�4  �|'  B� �q'  .��  �#/  )/  &8   /��  �:/  E/  &8  
8   0*  ���  �.  ^/  d/  ,8   0Ư  �p�  /  }/  �/  ,8   0�F  �5�  28  �/  �/  &8   0�F  �÷  �.  �/  �/  &8  
�2   0a�  ��j  28  �/  �/  &8   0a�   �i  �.  �/  	0  &8  
�2   0�:  m�  �.  "0  -0  ,8  
�.   0�F  	�u  28  F0  Q0  &8  
�.   0(*  �  �.  j0  u0  ,8  
�.   0 I  *�  28  �0  �0  &8  
�.   0�O  �  �.  �0  �0  ,8  
�.   0WC  �i  8  �0  �0  ,8    {�  �5   �  �   S�&  �,  �.  CU  A�7  1  
t8  
�2   D��  I01  
t8  
�2   D��  \F1  
t8  
�2   4Rj ��2  d1   �  �,  
�,   C9+  N�7  ~1  
t8  
�2   3�y  ��,  �1   {�  M5   �  �  
@B  
@B   3�v /�2  �1   {�  M5   �  �  
@B  
@B   3�l =�2  2   {�  M5   �  �  
@B  
@B   4;% ��2  #2   �   3  
M5   4��  ��2  A2   �  �5  
�5   3@k ��.  n2   {�  �5   �  �  
K  
K   #m /�r �2   {�  �5   �  �  
K  
K    E�  Eo  E�  E�  E�  E�  E�	  Fint E(  E#  E�� E�� E�� �2  E�  �2  2*  73  G8�    H�  E�  �  �2  �  �2  �O �2  �O �2  pW   �2  qW  !�2    "�2    #�2  ` &�2  ` '�2  �^ (�2  �^ )�2  �T *�2  �T +�2  iY ,�2  hY -�2  �e 0�2  �e 1�2  [ 2�2  [ 3�2  Q 4�2  Q 5�2  �_ 6�2  �_ 7�2  �] :�2  �] ;�2  �Q >�2  �Q ?�2  .  <^3  `  D�2  �  W^3  �  _i3  �  e�2  t   m�2  a  u�2    ~�2  �  ��2  3  ��2  �  ��2  H  ��2  y  ��2    ��2  s  ��2  T   ��2  �  ��2  F  ��2  �  ��2  �  ��2    ��2  V  ��2  I 3  E�  Js  N'3  �  V'3  \	  2�2  o  7�2  �  <�2  �  C�2  �  �2  I�5  KI�5   3  LpO qO !�5  M�   M�   I�   I�   M�  EYe E�[ I1  I�  M�  N1  M1  I�  M 3  M�5  IQ+  M�,  I�,  I�  M�  E  �  8|7  �{  M5   ]�  M5  \�   M5  �D  !M5  �3  "M5  U>  #M5  &�  $M5  �  %M5  �*  &M5   ڡ  ' 3  $�U  ( 3  %TL  ) 3  &�I  * 3  'Q  + 3  (�C  , 3  )�J  - 3  *1  .M5  ,o(  / 3  0�U  0 3  1PL  1 3  2�I  2 3  3Q  3 3  4�C  4 3  5�J  5 3  6 4)%  KM5  �7  
�2  
�5   OGT  P�7  IO6  �    �2  �2  I�  I�%  I�  I�  M�  M�%  N�  M�  P�2  �7  Q I�  I�,  M8  M5  I�0  M�,  IJ'  M!8  �5  I�.  I�0  M�.  I�%  I�'  Iz#  M%(  I%(  Mz#  IG!  M�(  I�(  MG!  I�7  R 1  �8  SXF  At8  S\;  A�2  TU�T  C�7    R1  �8  SXF  It8  S\;  I�2   R�   �8  ShR  ��8  SmR  ��8   �5  �5  R�   9  ShR  �9  SmR  �9   �5  �5  RH  N9  V__s 
�5  V__n 
W  V__a 
N9   �5  W�  !�Z5  t9  
W  X__p !�Z5   Y�  �9  �9  Zh  �9   �7  R�  �9  [�e  �5  [�e  �5  V__n W   Rl  �9  [�e  �5  [�e  �5  V__n W   R�  :  V__s �5  V__n W  V__a �    R
  M:  V__d dM5  V__s d�5  V__n d@   Y�  [:  e:  Zh  �9   Y�  s:  }:  Zh  �9   Y*  �:  �:  Zh  �9   Y"  �:  �:  Zh  �9  [%  D@   Yp	  �:  �:  Zh  �9  [%  A@  V__s A�5   Y�	  �:  ';  Zh  �9  [%  S@  [Q  S@  T\�c  U�2    R
  V;  [�e  �5  [�e  �5  V__n W   Y�  d;  n;  Zh  �9   R.  �;  V__s �5   R:  �;  T]__p �Z5    Y�  �;  �;  Zh  �;   �7  Y�  �;  �;  Zh  �;   Y�  �;  �;  Zh  �;  X__n �@   R01  <  SXF  \t8  S\;  \�2   YM&  $<  .<  Zh  .<   >8  Y/&  A<  K<  Zh  .<   Y
-  Y<  o<  Zh  o<  V__i �t<   �7  �7  Y'  �<  �<  Zh  �<  V__x n�<  V__y n�<   8  8  8  Y�.  �<  �<  Zh  �<   	8  R�
  =  V__p �M5  [۶  �M5  [nh  �M5   Y�0  =  =  Zh  =   ,8  R�
  P=  V__p �M5  [۶  ��5  [nh  ��5   Y)/  ^=  t=  Zh  t=  V__i �y=   &8  8  I�'  ^�'  v�=  �=  Zh  �=   ~=  Ia(  ^m(  v�=  �=  Zh  �=   �=  Y�  �=  �=  Zh  �9   Y�!  �=  >  Zh  >  X__x g!   \8  Y�  >   >  Zh  �9   R�(  >>  ;_Tp  3  
>>  
C>   B6  B6  M3  R�(  x>  ;_Tp �2  X__a �x>  X__b �}>   H>  H>  R�
  �>  [7i �@  [<i �@  T___d �    YS,  �>  �>  Zh  �>  X__p mi+  
]+   *6  RF1  �>   �  �,  
�,   Y�+  ?  ?  Zh  �>  Z#  �7   Ys  (?  ;?  Zh  ;?  Z#  �7   <6  Y�+  N?  ]?  Zh  �>  
]?   06  YX  p?  �?  Zh  ;?  X__a s�?   B6  Rd1  �?  SXF  Nt8  S\;  N�2   Y;  �?  �?  Zh  �;  X__a ��?   B6  Y�  �?  �?  Zh  �9   `  �?  @  Zh  @  Z#  �7   �7  M  `+  +@  :@  Zh  @  
:@   @  aN  Y�  S@  i@  Zh  i@  V__p (M5   �7  Y�+  |@  �@  Zh  �>   YB  �@  �@  Zh  ;?   Y�  �@  �@  Zh  @  [v�  M5  V__a �@   B6  Yw,  �@  �@  Zh  �@   66  Y+,  �@  A  Zh  �>  X__n c]+  
�5   Y�  &A  0A  Zh  �9   Yf  >A  HA  Zh  HA   �7  R,
  |A  V__d mM5  V__s m�5  V__n m@   Y�  �A  �A  Zh  �;   YI  �A  �A  Zh  HA   YV	  �A  �A  Zh  i@   Yx  �A  �A  Zh  i@   Y�#  �A  �A  Zh  �A  X__x �#   D8  YF  B  (B  Zh  i@  [%  U@   Y	  6B  @B  Zh  �9   M�0  R~1  {B   {�  M5   �  �  [\C  �{B  [?)  ��B   @B  @B  Y�	  �B  �B  Zh  �9  [7i K@  [<i K@  V__s K�5   RL
  �B  V__d vM5  V__n v@  V__c v 3   `x  �C  ;C  Zh  i@  [�m �@  [7i �@  [<i �@  V__c � 3   Y�  IC  kC  Zh  i@  V__n �@  V__c � 3   YK  yC  �C  Zh  i@  [��  Q�  [�  Q�  V__n Q@  V__c Q 3   `�  ��C  �C  Zh  i@  [�m �@  [7i �@  V__s ��5  [<i �@   Y�	  D  "D  Zh  �9  V__s [�5   b   �`D  V__n �@  V__c � 3  V__a �`D  T]__r ��7    B6  `  )vD  �D  Zh  i@  V__s ��5  V__n �@  T\R'  0Y  T\Q  7Y     `[  �D  �D  Zh  i@  V__n @  V__c  3  T\R'  Y    Y^  E  E  Zh  i@   Y�  E  .E  Zh  i@  Z#  �7   Yx  <E  FE  Zh  �;   Y�  TE  tE  Zh  �;  S�s �tE  S�s �yE   B6  B6  R�(  �E   8�  �,  
�E   @B  R)  �E   ��  �,  Sz  Z�,  S�l  Z�,  
n    R�1  F   {�  M5   �  �  [\C  /F  [?)  0F   {�  M5   �  �   @B  @B  R�1  QF   {�  M5   �  �  [\C  =QF  [?)  >VF   @B  @B  R?)  �F   f�  �,  Sz  r�,  S�l  r�,   Rl
  �F  V__p �M5  [۶  ��  [nh  ��   R  �F   �  �,  [�|  ��,  [�h  ��,  V__a ��F  
0   c B6  R:  0G   �  �,  [�|  ��,  [�h  ��,  V__a �0G  c B6  Y8	  CG  MG  Zh  �9   Y�  [G  qG  Zh  i@  [�^  *qG   �7  Rb)  �G   8�  M5  
�G   �7  R�)  �G   ��  M5  Sz  ZM5  S�l  ZM5  
n    R2  �G   �   3  SŐ  �M5   R�)  H   f�  M5  Sz  rM5  S�l  rM5   Rc  kH   ß  M5  S�|  |M5  S�h  |M5  X__a |kH  
H   daH  U�  �Y  ]__r ��7    ß  M5   B6  R�  �H   �  M5  [�|  �M5  [�h  �M5  V__a ��H  
0   c B6  R�  �H   �  M5  [�|  �M5  [�h  �M5  V__a ��H  c B6  R�)  
I   8�  �5  

I   8  R�)  >I   ��  �5  Sz  Z�5  S�l  Z�5  
n    R#2  ]I   �  �5  SŐ  ��5   R*  �I   f�  �5  Sz  r�5  S�l  r�5   R�  �I   ß  �5  S�|  |�5  S�h  |�5  X__a |�I  
H   d�I  U�  �Y  ]__r ��7    ß  �5   B6  R   )J   �  �5  [�|  ��5  [�h  ��5  V__a �)J  
0   c B6  RB   gJ   �  �5  [�|  ��5  [�h  ��5  V__a �gJ  c B6  Y�  zJ  �J  Zh  i@  [��  '�  [�  '�  V__s '�5  V__n '@   Yk&  �J  �J  Zh  .<   Y�  �J  K  Zh  i@  [��  ��  [�  ��  [۶  ��5  [nh  ��5   M�0  RA2  OK   {�  �5   �  �  [\C  �OK  [?)  �TK   K  K  et9  n%  p|   �tK  }K  f�9  �  eE@  �I  �|   ��K  �K  fS@  � f\@  � eM:  �%  �|
   ��K  �K  f[:  �  e(B  E)  �|   ��K  L  f6B  �gK<  �|`�  3hb<  fY<  �   e5G  ;&  �|   �*L  nL  fCG  �it9  �|x�  7OL  f�9  � jK<  �|   7hb<  fY<  �   e�:  :2  �|(   ��L  �L  f�:  � f�:  �f�:  �ie:  �|��  C�L  fs:  �  k�|�*   e�B  �(   }+   ��L  *M  f�B  � f�B  �f�B  �f�B  �le:  }   M M  fs:  �  k+}
+   e�:  >$  0}   �EM  �M  f�:  � f ;  �f;  �m��  n;  � <�@K$"�@K$"+�ge:  0}��  Ufs:  �    e�C  �7  P}   ��M  �M  fD  � fD  �gt9  P}��  ]f�9  �   o:  �-  p}6   �kN  p(:  � p4:  >� p@:  h� l�9  �}"   iKN  p�9  �� p�9  �� p�9  ܨ q�}�   j�8  �}   gf�8  Qf�8  R  oMA  �P  �}6   ��N  pWA  �� pcA  %� poA  O� l�9  �}"   r�N  p�9  �� p�9  �� p�9  é q�} �   j�8  �}   pf�8  Qf�8  R  o�B  \-  �}3   ��O  p�B  � p�B  � p�B  6� l�9  ~   {aO  p:  V� p:  i� p�9  �� q~B�   j�8   ~   yf�8  �  f�8  Q  o�F  �-  0~6   �fP  p�F  �� p�F  Ѫ f�F  �g�<  4~��  �p�<  �� p�<  &� p�<  F� j:  >~(   �p@:  p� p4:  �� p(:  �� l�9  C~    iFP  p�9  � p�9  �� p�9  � qT~�   j�8  c~   gh�8  f�8  Q    r�
  p~6   �WQ  s__p �M5  0� t۶  ��  Z� unh  ��  �g!=  t~�  �pC=  �� p7=  �� p+=  Ϭ j:  ~~(   �p@:  �� p4:  )� p(:  I� l�9  �~    i7Q  p�9  s� p�9  �� p�9  �� q�~�   j�8  �~   gh�8  f�8  Q    o�<  �   �~6   �R  p�<  �� p�<  � p�<  � j:  �~(   �p@:  -� p4:  \� p(:  �� l�9  �~    i�Q  p�9  �� p�9  î p�9  � q�~�   j�8  �~   gh�8  f�8  Q   o!=  IP  �~6   ��R  p+=  � p7=  +� pC=  U� j:  �~(   �p@:  u� p4:  �� p(:  ί l�9      i�R  p�9  �� p�9  � p�9  *� q�   j�8  #   gh�8  f�8  Q   o�>  rR  0	   ��R  f�>  � f�>  �v0   w�>  I�   x?@  D*  @   �e�D  �p P   �*S  ZS  fE  � j�@  P   �h�@  p�@  n� f�@  �   Yk  hS  ~S  Zh  i@  [�^   ~S   �7  eZS  Dw `   ��S  �S  fhS  � fqS  �l@  d   �S  f4@  �f+@  �  jE@  l   p\@  �� fS@  �  e>  �>  �   �T  8T  f>  �gP=  � �  rhg=  f^=  �   e�=  6;  �   �ST  �T  f�=  �it9  �8�  �xT  f�9  � jP=  �   �hg=  f^=  �   y  �   ��T  U  zh  �9  �i�=  �P�  ��T  f�=  �gt9  �h�  �f�9  �  j�=  �   �p�=  �� f�=  �   yQ  �   �*U  YU  zh  �9  �g�=  ���  �p�=  � f�=  �   yp  �   �pU  �U  zh  �9  �gP=  ���  �hg=  f^=  �   y�  �   ��U  �U  zh  �9  �it9  ���  ��U  f�9  � jP=  �   �hg=  f^=  �   y�  �   �V  vV  zh  �9  �i�=  ���  �SV  f�=  �gt9  ���  �f�9  �  j�=  �   �p�=  � f�=  �   y�  0�   ��V  �V  zh  �9  �g�=  0���  �p�=  ,� f�=  �   ee:  �R  @�
   ��V  �V  fs:  �  y  P�
   ��V  W  zh  �9  �  e}:  j=  `�   �W  (W  f�:  �  eA  v  p�
   �CW  LW  f&A  �  y  ��   �cW  �W  zh  �9  � je:  ��   6fs:  �   e�:  �6  ��   ��W  �W  f�:  � f�:  � yj  ��'   ��W  @X  zh  �9  � {__n k@  �ie:  ���  m6X  fs:  � gM:  ��(�  �f[:  � gt9  ��(�  -f�9  �    kǀ�*   y�  Ѐ   �WX  dX  zh  �9  �  y  ��   �{X  �X  zh  �9  � le:  ��   ��X  fs:  � jM:  ��   �f[:  � jt9  ��   -f�9  �    j�:  �   �p�:  P� f�:  �   |$  ���q   �Y  �Z  zh  �9  � {__s M5  �s__n @  u� u%  @  �i�:  �@�  ��Y  f�:  �	�p�:  �� f�:  � ie:  �`�  C�Y  fs:  � gM:  �x�  �f[:  � gt9  �x�  -f�9  �    ka��*   l�:  	�   �Z  p;  ˱ p ;  � p�:   � v	�   w;  4�   g:  ���  �p@:  ˲ p4:  �� p(:  #� l�9  �   i~Z  p�9  C� p�9  V� p�9  i� k)��   j�8  C�   gh�8  p�8  }�    |R  p�9   ��Z  �[  }h  i@  �� s__s �[  �� lM:  y�   	[  p[:  ϳ jt9  y�   -p�9  ϳ   lM:  ��   F[  p[:  � jt9  ��   -p�9  �   l�;  ��   d[  p�;  �  ~��   �[  \Y�  M5  lE@  ��   �[  p\@  � pS@  *�  jE@  ��   p\@  >� pS@  Q�   j�;  ��	   
f�;  rt�  �7  y0  ��   ��[  $\  zh  i@  � u�^  M$\  �k�Z   �7  y�  Ё   �@\  e\  zh  i@  � u�^  Ie\  �k��Z   �7  yr  ��   ��\  �\  zh  �9  �  eV;  �A   �   ��\  �\  fd;  �  e�?  Z5  �   ��\  �\  f�?  � |�  � ��   ��\  �]  zh  �9  � {__s <�5  �t%  <@  e� {__n <@  �m��  \�a  �Y  \�k ��5  ie:  '���  ��]  ps:  ʴ gM:  '���  �p[:  ʴ gt9  '���  -p�9  ʴ    j';  ��   �pI;  �� p=;  � p1;  E� k��d�     y�  ��   ��]  j^  zh  �9  � u�^  Ij^  �u%  I@  �le:  �   K`^  fs:  �jM:  �   �f[:  �jt9  �   -f�9  �   k
��\   �7  y&  �%   ��^  �^  zh  �9  � {__s X�5  �u%  X@  �ln;  �	   [�^  px;  c� k���   k0��\   |O  �@�T   ��^  `  zh  �9  � {__c i 3  �u%  i@  �m �  �&  �@  �� \�a  �Y  ie:  C� �  ��_  fs:  � gM:  C�8�  �f[:  � gt9  C�8�  -f�9  �    vp�   \�k ��5  �__n �Y  е ___p  �5  g9  p�P�   fA9  �*6  p59  е p)9  �� k����      |�  	��}   �`  �`  zh  �9  � {__s ��5  �t%  �@  )� {__n �@  �mx�  \�a  Y  ie:  ����  �`  fs:  � gM:  ����  �f[:  � gt9  ����  -f�9  �    m��  \�k �5  j';  �   pI;  v� p=;  �� p1;  � k��d�      yx   �   �a  �a  zh  �9  � u�^  v�a  �u%  v@  �le:  #�   x�a  fs:  �jM:  #�   �f[:  �jt9  #�   -f�9  �   k:�`   �7  y�  @�%   ��a  b  zh  �9  � {__s ��5  �u%  �@  �ln;  H�	   �b  px;  5� kN���   k`�`   |�  p�A   �*b  �b  zh  �9  � s__c � 3  T� u%  �@  �m��  �a  !@  � ge:  q��  !fs:  � gM:  q�8�  �f[:  � gt9  q�8�  -f�9  �      |J  /��j   ��b  �c  zh  �9  � {__s ��5  �t%  �@  �� {__n �@  �le:  ؄	   3]c  ps:  ҷ jM:  ؄   �p[:  ҷ jt9  ؄   -p�9  ҷ    mP�  ___p 5�5  j9  ��   5pA9  � p59  <� p)9  f� k���     y!  0�   ��c  ?d  zh  �9  � u�^  �?d  �u%  �@  �le:  3�   �5d  fs:  �jM:  3�   �f[:  �jt9  3�   -f�9  �   kJ��b   �7  yx  P�%   �[d  �d  zh  �9  � {__s ��5  �u%  �@  �ln;  X�	   ��d  px;  �� k^���   kp��b   y�  ��   ��d  e  zh  �9  � s__c � 3  �� u%  �@  �����^  �� � ���  |�  >��i   �0e  f  zh  �9  � {__s �5  �u%  @  �{__n @  �mh�  �a  B@  ĸ ie:  ����  B�e  ps:  � gM:  ����  �p[:  � gt9  ����  -p�9  �    j9  م   IpA9  >� p59  f� p)9  �� k���     y�   �   �f  �f  zh  �9  � u�^  ��f  �u%  �@  �le:  �   ��f  fs:  �jM:  �   �f[:  �jt9  �   -f�9  �   k�e   �7  y!   �%   ��f  g  zh  �9  � {__s �5  �u%  @  �ln;  (�	   g  px;  �� k.���   k@�e   yJ  P�   �/g  xg  zh  �9  � s__c $ 3  ù u%  $@  ��^�b  �� � ���  |�  S`�m   ��g  Th  zh  �9  � {__s C�5  �t%  C@  � {__n D@  �ie:  g���  Wh  ps:  � gM:  g���  �p[:  � gt9  g���  -p�9  �    j9  ��   XpA9  6� p59  p� p)9  �� k����    ys  І   �kh  �h  zh  �9  � u�^  2�h  �u%  2@  �le:  ӆ   4�h  fs:  �jM:  ӆ   �f[:  �jt9  ӆ   -f�9  �   k�xg   �7  y�  ��%   �
i  ei  zh  �9  � {__s Q�5  �u%  Q@  �ln;  ��	   T[i  px;  �� k����   k�xg   |�  _ �E   �i  �i  zh  �9  � {__c b 3  �t%  b@  ͺ ge:  #��  bfs:  � gM:  #� �  �f[:  � gt9  #� �  -f�9  �     |E  jp�}   �j  �j  zh  �9  � {__s ��5  �u%  �@  �{__n �@  �m8�  �a  n@  � ie:  w�h�  n�j  fs:  � gM:  w���  �f[:  � gt9  w���  -f�9  �    j9  ��   upA9  H� p59  �� p)9  �� kȇ��     y  ��   ��j  ~k  zh  �9  � u�^  q~k  �u%  q@  �le:  �   stk  fs:  �jM:  �   �f[:  �jt9  �   -f�9  �   k
��i   �7  ys  �%   ��k  �k  zh  �9  � {__s ��5  �u%  �@  �ln;  �	   ��k  px;  � k���   k0��i   |�  @�G   �l  �l  zh  �9  � s__c � 3  � u%  �@  �m��  �a  �@  6� ge:  A���  �fs:  � gM:  A���  �f[:  � gt9  A���  -f�9  �      y�  ��3   ��l  n  zh  �9  � u�^  �n  �v��(   �a  �Y  �� /i �Y  �� \R'  �Y  �__r ��2  Pie:  ����  �am  fs:  � gM:  ���  �f[:  � gt9  ���  -f�9  �    ie:  ��0�  ��m  fs:  �gM:  ��P�  �f[:  �gt9  ��P�  -f�9  �   i�>  ��h�  ��m  h�>  h�>  mh�  ��>    j';  ��   �hI;  p=;  �� p1;  Ǽ k��d�     �7  |  �Ј[   �-n  p  zh  �9  � t%  �@  ڼ s__n �@  � u�^  �p  �m��  /i �Y  p� \R'  �Y  �__r ��2  �� i�:  ӈ��  �$o  f�:  �	�p�:  �� f�:  � ie:  ӈ��  Co  fs:  � gM:  ӈ��  �f[:  � gt9  ӈ��  -f�9  �    k+��*   l�:  �   �go  p;  �� p ;  ս p�:  � v�   w;  ��   ie:  ���  ��o  ps:  b� gM:  ��  �p[:  b� gt9  ��  -p�9  b�    i';  � �  ��o  hI;  p=;  v� p1;  �� k�d�   g�>  �8�  �h�>  h�>  m8�  ��>      �7  |@  �0��   �6p  �r  zh  �9  � u�m �@  �t7i �@  �� u�^  ��r  �u�m �@  �t<i �@  ؾ mP�  \R'  �Y  �__r ��2  � i�:  7�p�  �?q  f�:  �	�p�:  "� p�:  o� ie:  7���  C5q  ps:  o� gM:  7���  �p[:  o� gt9  7���  -p�9  o�    k���*   i�:  P���  ��q  p�:  �� p�:  Ϳ p�:  �� le:  P�	   C�q  ps:  �� jM:  P�   �p[:  �� jt9  P�   -p�9  ��    k���*   l�:  ]�   �r  p;  � p ;  6� p�:  U� v]�   w;  i�   l�:  d�   �Pr  p;  �� p ;  �� p�:  � vd�   w;  *�   i';  o���  ��r  hI;  p=;  �� p1;  �� k��d�   j�>  ��   �h�>  h�>  v��   ��>      �7  |x  ���=   ��r   t  zh  �9  � {__s 	�5  �m��  �a  �Y  �� /i �Y  � \R'  �Y  �__r ��2  Pie:  ǉ�  �{s  fs:  � gM:  ǉ �  �f[:  � gt9  ǉ �  -f�9  �    ln;  ԉ   ��s  px;  "� kډ��   i�>  �8�  ��s  h�>  h�>  m8�  ��>    j';  �   �hI;  p=;  A� p1;  `� k��d�     |�  � �j   �t  �u  zh  �9  � u%  (	@  �t7i (	@  s� {__s (	�5  �mP�  /i �Y  �� \R'  �Y  �__r ��2  �� i�:  �p�  �u  f�:  �	�p�:  �� p�:  �� ie:  ���  C
u  ps:  $� gM:  ���  �p[:  $� gt9  ���  -p�9  $�    kj��*   l�:  �   �Wu  p;  O� p ;  n� p�:  �� v�   w;  ��   ln;  #�   �~u  px;  �� k/���   i�>  ?���  ��u  h�>  h�>  m��  ��>    j';  A�   �hI;  p=;  �� p1;  � kL�d�     |�  �p�Z   ��u  �w  zh  �9  � u%  C	@  �t7i C	@  L� {__s C	�5  �u<i D	@  �m��  \R'  �Y  �__r ��2  �� i�:  u���  ��v  f�:  �	�p�:  �� f�:  � ie:  u��  C�v  fs:  � gM:  u�0�  �f[:  � gt9  u�0�  -f�9  �    kʊ�*   l�:  ��   �.w  p;  �� p ;  � p�:  1� v��   w;  E�   i';  ��H�  �cw  hI;  p=;  �� p1;  �� k��d�   g�>  ��`�  �h�>  h�>  m`�  ��>      e�@  Np Њ   ��w  �w  f�@  � f�@  �f�@  � x�;  �O  ��   �e�A  �N  ��   ��w  �w  f�A  �  e0A  o+   �   �x  x  f>A  �  e|A  �O  �   �6x  ?x  f�A  �  e�;  �P   �   �Zx  cx  f�;  �  e�;  -  0�#   �~x  �x  f�;  � f�;  �v@�   f�;  �f�;  � ��;  D�   ��x  f�;  �  ��8  M�   �h�8  f�8  
� �"#�   e�;  �R  `�   �y  y  f�;  �  r  p�v   �.z  t� "@  �� u�t "@  �u�o #.z  �mx�  $t AY  I� +k BY  _� �a  P@  s� zs RY  �� <w _Z5  � ___p `�7  ~��   �y  �p UY  +�  l�@  ��	   _z  h�@  pA  �� pA  �� kʋ��   l�;  ͋   i#z  p�;  ��  k�
+    B6  o"D  3J  ���   ��{  f.D  � f:D  �fFD  ����  sz  �SD   m��  pFD  �� p:D  �� p.D  � m��  wSD  =� ��B  ���  �-{  p�B  q� p�B  �� p�B  �� l�9  $�   {	{  p:  �� p:  
� p�9  � k4�B�   j�8  P�   yp�8  0� p�8  H�   ��;  �   �K{  p�;  =�  ��;  7���  ��{  p�;  [� p�;  y� v`�   f�;  Sf�;  W��;  `�   դ{  f�;  W ��8  i�   �h�8  f�8  w s "#�   k�y     ^u  � �{  �{  Zh  i@  V__a ��{   B6  e�{  �w p�   �|  b|  f�{  � f�{  ���@  ��   �X|  f�@  �f�@  Pf�@  �  k��"D   ^E  � r|  �|  Zh  i@  V__n �@  V__c � 3  V__a ��|   B6  eb|  �v ��    ��|  }  fr|  � f{|  �f�|  �f�|  ���@  ��   �}  f�@  �f�@  Pf�@  �  k��"D   r�  ��   �u}  u�i �@  � s__c � 3  �� {__a �u}  ����"D  �� � ���  B6  yY  ��   ��}  ~  zh  �;  � {__a �~  �v��   �a  �Y  �� j�>  ��   �h�>  p�>  �� f�>  � �Ō��  �� �     B6  ��?  Ќ2   �~  �~  p�?  �� p�?  �� ��?  Ԍ��  ��~  ��?  p�?  � �z8  Ԍ��  V��8  p�8  � m��  w�8  8�    k��z}   e�?  |6  �#   ��~  3  f�?  � f�?  �m�  h�?  f�?  � ��?   �(�  �(  ��?  f�?  � #��z8   �(�  V��8  f�8  � #�m(�  w�8  X�    q3�z}    eE  x @�@   �N  *�  fE  � lM:  D�	   #�  f[:  � jt9  D�   -f�9  �   g�?  M�@�  #p�?  k� p�?  �� v`�    p�?  �� p�?  �� ��?  `�X�  ��  ��?  p�?  �� �z8  `�X�  V��8  p�8  �� mX�  w�8  �    k{�z}     |  ����  �D�  ��  zh  i@  � u%  �@  �u�m �@  �u�m �@  �mp�  \�t �Y  ]8 �Y  +� gr �Y  T� ie:  ����  ���  fs:  � gM:  ����  �f[:  � gt9  ����  -f�9  �    lA  ��   ��  f&A  �  ���  ��  �__a �k   �_�__r ��7  }� it9  ύ��  �c�  p�9  ��  i:  Ӎ�  ��  p@:  �� p4:  � p(:  1� l�8  �   g��  h�8  p�8  [�  j�9  �   ip�9  n� p�9  �� p�9  �� k��    i�;  ֍0�  �	�  p�;  ��  lM:  ��	   �A�  p[:  �� jt9  ��   -p�9  ��   i�?  �H�  �ނ  p�?  �� p�?  (� v �#   f�?  Sp�?  F� ��?   �`�  �ӂ  ��?  p�?  Y� �z8   �`�  V��8  p�8  Y� m`�  n�8  V   k;�z}    iE@  �x�  ��  p\@  n� pS@  ��  i:  F���  ���  p@:  �� p4:  �� p(:  �� l�8  R�   gW�  h�8  p�8  �  j�9   �    ip�9  � p�9  -� p�9  @� k��    kƍy   iMA  |���  ��  poA  S� pcA  q� pWA  �� l�8  ��   p�  h�8  p�8  ��  j�9  ��$   rp�9  �� p�9  �� p�9  �� kˎ �    g�;  ���  �p�;  � p�;  .� v��   p�;  P� h�;  ��;  ��   �r�  h�;   ��8  ��   �h�8  p�8  c�      |4  �P�5   ���  �  zh  i@  � lM:  X�   ��  f[:  � jt9  X�   -f�9  �   l|A  y�   ��  p�A  {�  kt�*�   e�A  �>  ��"   �4�  o�  f�A  � l�A  ��   <Z�  p�A  ��  �����  �� �   e�A  �&  ��0   ���  �  f�A  �l�A  ͏   h�  p�A  �� lM:  ͏   <�  p[:  �� jt9  ͏   -p�9  ��   kߏ��   jK<  �   ihb<  pY<  ��   y2  ��0   �(�  ц  zh  i@  �l�A  ��   ���  p�A  �� j�A  ��   hp�A  �� lM:  ��   <��  p[:  �� jt9  ��   -p�9  ��   k���    j�A  �   �f�A  R�p�A  �   Y�  ߆  �  Zh  i@   eц  <   �3   ��  ��  f߆  �l�A  -�   {k�  p�A  0� lM:  -�   <a�  p[:  0� jt9  -�   -p�9  0�   k?���   jK<  I�   |hb<  pY<  O�   eB  W  `�(   ���  �  fB  � fB  �j�A  h�   \f�A  � lM:  h�   <�  f[:  � jt9  h�   -f�9  �   kz���    y�  ��$   �&�  ��  zh  i@  � jB  ��   ��B   fB  � j�A  ��   \f�A  � lM:  ��   <��  f[:  � jt9  ��   -f�9  �   k����     y�  ��.   �  b�  zh  i@  � le:  ɐ   ��  fs:  � jM:  ɐ   �f[:  � jt9  ɐ   -f�9  �    gB  ѐ��  �pB  m� fB  � j�A  ѐ   \f�A  � k���     y�  �@   �y�  �  zh  i@  � {__n �@  �le:  ��   ��  ps:  �� jM:  ��   �p[:  �� jt9  ��   -p�9  ��    l�A  �   ��  p�A  �� k���   k0��*   y�  0�3   �.�  ׊  zh  i@  �lц  =�   ���  p߆  �� j�A  =�   {p�A  �� lM:  =�   <��  p[:  �� jt9  =�   -p�9  ��   kO���    j�A  Y�   �p�A  �� p�A  ��   y�  p�   ��  "�  zh  i@  � le:  y�   .�  ps:  �  k��*�   Y1  0�  R�  Zh  i@  [%  d@  V__n d@   e"�  �R  ��F   �m�  (�  f0�  � f9�  �fE�  �l�:  ��   g�  p;  7� p ;  a� p�:  �� v��   w;  �� je:  ��   Ups:  ��    i�:  ����  g�  f�:  F��p�:  � p�:  I� k֑�*   k��*�   yZ  ��4   �?�  ��  zh  i@  �tv t�  h� m�  %  xY  �� iFB  �(�  x��  hnB  fbB  �nc   lM:  ��   z̌  f[:  �jt9  ��   -f�9  �  l|A  �   z�  p�A  ��  k��*�    |~  � �X   ��  �  zh  i@  �tz  ��  �� u�l  ��  �m@�  �a  �Y  �� vD�-   %  �Y  � lFB  D�   ���  hnB  fbB  �>d   lM:  Y�   �č  f[:  �jt9  Y�   -f�9  �  lK<  c�   ��  hb<  hY<   l|A  f�   ��  p�A  (�  kY�*�     e�B  �&  ���   �(�  }�  fC  � f
C  �fC  �f"C  �f.C  �i�B  ��`�  ���  f�B  �	�p�B  N� p�B  �� p�B  �� le:  ��	   M��  ps:  ��  k�
+   �x�  s�  pC  � p.C  &� p"C  Z� p
C  �� pC  �� g�B  ����  �p�B  �� p�B  � p�B  7� l�9  Œ   {N�  p:  U� p:  ~� p�9  �� kՒB�   j�8  �   yp�8  �� p�8  ��    k��*�   e;C   @  �"   ���  ؏  fIC  � fRC  �f^C  �le:  !�   �Ώ  ps:  ��  k.��B   y  @�$   ��  [�  zh  i@  � {__c = 3  �g;C  D���  ?f^C  ��RC  pIC  �� le:  N�   �P�  ps:  ��  k]��B    y�  p�A   �r�  �  zh  i@  � u%  9@  �{__n 9@  �{__c 9 3  �i�:  ����  ;�  f�:  	�p�:  � p�:  B� le:  ��   C��  ps:  B�  k���*   k���B   y  ��=   �&�  �  zh  i@  �s__p K�  x� {__c K 3  �m��  %  NY  �� iFB  ˓��  N��  hnB  fbB  �Uh   lM:  �   P  f[:  �jt9  �   -f�9  �  l|A  �   P��  p�A  ��  k��B    y�   �_   ��  �  }h  i@  �� t%  @  �� t7i @  � t<i @  0� s__c  3  P� l�:  �   ��  p;  p� p ;  �� p�:  �� v�   w;  �� je:  �   Ups:  ��    i�:  *��  �  f�:  	�p�:   � p�:  J� k_��*   qN��B   ekC  'S  `�&   ��  ��  fyC  � p�C  t� f�C  �f�C  �p�C  �� lFB  q�   Ud�  fnB  �  fbB  �   lFB  {�   U��  hnB  fbB  �   ����B  �� � ���  y�  ��$   ���  g�  zh  i@  � s__p ��  �� {__n �@  �{__c � 3  �gkC  �� �  �f�C  �f�C  �f�C  ��f�C  ��pyC  �� lFB  ��   U\�  hnB  fbB  �Fk   k���B    e�C  O  ��O   ���  p�  f�C  � f�C  �f�C  �f�C  �f�C  ��8�  f�  p�C  �� p�C  � p�C  G� p�C  g� p�C  �� g:  �P�  �p@:  �� p4:  �� p(:  �� l�9  �   iE�  p�9  � p�9  /� p�9  C� k���   j�8  �   gh�8  p�8  V�    k۔*�   |>  ��   ���  �  }h  i@  i� s__s n�5  �� s__n n@  � ie:  �h�  	�  ps:  .� jM:  �   �p[:  .� jt9  �   -p�9  .�    i�B  !���  N�  f�B  3	�p�B  z� p�B  �� p�B  �� kƕ
+   l�C  0�   u�  pD  I� pD  ��  ~W�b   ��  %  Y  �� l:  _�   ��  p@:  � p4:  *� p(:  I� j�9  d�   ip�9  \� p�9  o� p�9  �� ko��    l�;  t�   w�  p�;  �� p�;  �� v~�   p�;  �� p�;  �� ��;  ~�   �V�  p�;  ��  ��8  ��   �h�8  p�8  ��    jMA  ��%   poA  	� pcA  � pWA  ;� l�9  ��   rۗ  p�9  N� p�9  a� p�9  �� k�� �   j�8  ��   ph�8  p�8  ��    kI��C   yT  Е   ��  B�  zh  i@  � {__l Y�%  �k�p�   y  �L   �Y�  i�  }h  i@  �� t�^  ^i�  �� t%  ^@  �� s__n ^@  '� i�:  ���  a#�  p;  F� p ;  e� p�:  �� m��  w;  �� ge:  ���  Ups:  �� gM:  ���  �p[:  �� gt9  ���  -p�9  ��      i�:  ���  `_�  f�:  3	�p�:  �� p�:  � k<��*   q+�p�   �7  Yg  |�  ��  Zh  i@  V__s z�5   en�  �T  @�!   ���  �  f|�  � f��  �ln;  H�	   }�  px;  ;� kN���   k\�p�   y�  p�   ��  5�  zh  i@  � {__l ��%  ��u�p�  �� �   y�  ��!   �L�  ��  zh  i@  � {__s 2�5  �jn�  ��   3p��  Z� f|�  � ln;  ��	   }��  px;  Z� k����   k��p�    |�  g��q  �Ԛ  ��  zh  i@  � u%  @  �s__s �5  y� {__n @  �i�:  ǖ �  k��  f�:  	�p�:  �� p�:  *� le:  ǖ   C��  ps:  �� jM:  ǖ   �p[:  �� jt9  ǖ   -p�9  ��    k��*   i�B  Ԗ�  lޛ  p�B  �� p�B   � p�B  y� p�B  �� k!�
+   i�C  �0�  m�  pD  �� pD  U�  �H�  ��  Q  rY  �� �__p uM5  �� lt9  �   tN�  p�9  *�  i:  ,�p�  w֜  p@:  j� p4:  �� p(:  �� l�9  1�   i��  p�9  �� p�9  �� p�9  � k<��   g�8  ����  gh�8  p�8  �   ���  ��  �s |Y  (� i:  X���  }x�  p@:  (� p4:  F� p(:  d� l�8  d�   gB�  h�8  p�8  ��  j�9  �   ip�9  �� p�9  �� p�9  �� k���    g:  n���  ~p@:  �� p4:  � p(:  ,� l�8  v�
   gƝ  h�8  p�8  J�  j�9  З    ip�9  ]� p�9  �� p�9  �� kۗ�     i:  ����  y��  p@:  �� p4:  �� p(:  �� l�8  ��   gO�  h�8  p�8  �  j�9  ��    ip�9  $� p�9  7� p�9  J� k���    k�*�   k���C   y  0�   ���  �  zh  i@  � s__p ��  ]� {__l ��%  �lFB  4�   ��  hnB  fbB  ��u   �C���  �� �   YP  $�  ^�  Zh  i@  [�m �@  [�^  �^�  [�m �@  V__n �@   �7  e�  u>  P�\   �~�  }�  p$�  |� p-�  �� p9�  �� pE�  �� fQ�  �i�:  W��  �7�  p;  �� p ;  &� p�:  \� m�  w;  �� ge:  W� �  Ups:  \� gM:  W�8�  �p[:  \� gt9  W�8�  -p�9  \�      i�:  y�P�  �s�  f�:  	�p�:  �� p�:  � k���*   q����   y�  ��%   ���  �  zh  i@  � u%  "@  �{__s "�5  �ln;  ��	   %�  px;  7� k����   kИ��   y'  ��   ��  ¡  zh  i@  � u�m �@  �u�^  �¡  �le:  �   ��  fs:  �jM:  �   �f[:  �jt9  �   -f�9  �   j�  �   �pQ�  V� �E�   f9�  �f-�  �f$�  � k����    �7  y�   �3   �ޡ  x�  zh  i@  � le:  �   ��  ps:  ��  g"�  �h�  ��E�  p9�  �� p0�  �� i�:  ���  gm�  f�:  F��p�:  �� p�:  �� k3��*   k�*�    e.E  �-  @�   ���  ��  p<E  �� i�;  K���  ��  p�;  !�  j�;  P�   �
<  p�;  L� ��8  P�   d��8  p�8  L�    y�  `��   ��  ��  zh  �;  � u�o p��  �u/t  p@  �m��  �i sY  q� �__r t�7  �� i:  ����  w�  p@:  �� p4:  �� p(:  -� l�9  ��   i̣  p�9  a� p�9  t� p�9  �� k���   j�8  ʙ   gh�8  p�8  ��   i�;  ����  w
�  p�;  ��  l�;  ��   w(�  p�;  ��  i�;  ���  y��  p�;  � p�;  3� vә   f�;  Rp�;  k� ��;  ә   Յ�  p�;  k�  ��8  ܙ   �h�8  p�8  ��    k}�y    B6  |�  ���   �Ф  ��  zh  i@  � t/t  &@  �� lA  ��   �>�  p&A  � jM:  ��   p[:  � jt9  ��   -p�9  �    m(�  �__a �k   �_Y�  �M5  @� le:  �   ���  ps:  j�  lM:  �   ���  p[:  ��  iM:  "�@�  �ץ  p[:  �� jt9  "�   -p�9  ��   i�?  $�X�  �p�  h�?  p�?  �� vP�$   f�?  Vp�?  �� ��?  P�x�  �e�  ��?  p�?  �� �z8  P�x�  V��8  p�8  �� mx�  n�8  W   kk�z}    lE@  2�    ��  p\@  
� pS@  �  k"���    y�  ��B   ���  3�  zh  i@  � lA  ��   �  p&A  0� jM:  ��   p[:  0� jt9  ��   -p�9  0�    k����  k����  q�   |�  DК�   �M�  �  zh  i@  � u�^  ��  �m��  \�a  GY  le:  ߚ   G˧  ps:  s� jM:  ߚ   �p[:  s� jt9  ߚ   -p�9  s�    m��  R'  JY  �� le:  �   J2�  ps:  �� jM:  �   �p[:  �� jt9  �   -p�9  ��    i:  ���  M��  p@:  �� p4:  �� p(:  � l�9  �   i��  p�9  3� p�9  F� p�9  Y� k��   j�8  S�   gh�8  p�8  l�   lM:  �   N�  p[:  � jt9  �   -p�9  �   i�;   ���  Ns�  p�;  �� p�;  �� v`�   f�;  Uf�;  pt���;  `�   �O�  f�;  pt� ��8  j�   �h�8  f�8  p u "�   k����     �7  y,  p�   ���  ԩ  zh  i@  � u�^  �ԩ  ��u�3�  �� � ���  �7  |�  U���   ��  ��  zh  i@  � u�^  ���  �u%  �@  �s__n �@  �� i�:  ����  X��  f�:  H	�p�:  �� p�:  '� ie:  ��  C��  ps:  '� gM:  ��(  �p[:  '� gt9  ��(  -p�9  '�    kA��*   l�:  ��   Y��  p;  ]� p ;  |� p�:  �� v��   w;  ��   m@  R'  \Y  >� le:  ��   \e�  ps:  \� jM:  ��   �p[:  \� jt9  ��   -p�9  \�    i:  ؛X  _�  p@:  z� p4:  �� p(:  �� l�9  ݛ   iͫ  p�9  �� p�9  �� p�9  �� k��   j�8  �   gh�8  p�8  �   lM:  �   `%�  p[:   � jt9  �   -p�9   �   i�;  �p  `��  p�;  >� p�;  \� v �   p�;  ~� p�;  �� ��;   �   Մ�  p�;  ��  ��8  *�   �h�8  p�8  ��    kƛ��    �7  eeD  �D  P��   �Ь  [�  fvD  � fD  �f�D  �m�  p�D  �� pD  �� pvD  � m�  w�D  /� i�B  g��  /��  p�B  M� p�B  �� p�B  u� p�B  � ie:  g��  M��  ps:  � jM:  g�   �p[:  � jt9  g�   -p�9  �    k�
+   i�C  ���  3ѭ  pD  �� pD  ��  ~�   �  w�D  �� lt9  �   9�  p�9  �  k���   i:  ���  <��  p@:  � p4:  B� p(:  k� l�8  ��   ga�  h�8  p�8  ��  j�9  М   ip�9  �� p�9  �� p�9  �� kۜ�    lM:  ��   =Ϯ  p[:  �� jt9  ��   -p�9  ��   i�;  �� =O�  p�;  �� p�;  � v �   p�;  3� p�;  F� ��;   �   �.�  p�;  F�  ��8  
�   �h�8  p�8  [�    k����     y�   �   �r�  ��  zh  i@  � {__l ��%  ��%�eD  �� �   Y7  ��  Ư  Zh  i@  V__s ��5   e��  �*  0�!   ��  "�  f��  � f��  �ln;  8�	   �  px;  s� k>���   kL�eD   y�  `�   �9�  i�  zh  i@  � {__l �%  ��e�eD  �� �   yP  p�!   ���  �  zh  i@  � {__s ��5  �j��  x�   �p��  �� f��  � ln;  x�	   �  px;  �� k~���   k��eD    e�D  �6  ���   �	�  3�  f�D  � f�D  �f�D  �m  p�D  �� p�D  �� p�D  � m  w�D  ,� i�B  ��8 �  p�B  J� p�B  �� p�B  r� p�B  � ie:  ��P Mٱ  ps:  � jM:  ��   �p[:  � jt9  ��   -p�9  �    kM�
+   i�B  �h !o�  p�B  �� p�B  �� p�B  �� l�9  �   {K�  p:  � p:  +� p�9  >� k��B�   j�8   �   yp�8  Q� p�8  i�   lM:  ��   "��  p[:  |� jt9  ��   -p�9  |�   i�;  ��� "'�  p�;  �� p�;  �� v0�   p�;  �� p�;  �� ��;  0�   ��  p�;  ��  ��8  :�   �h�8  p�8  �    kٝ��     |I  P�w   �M�  u�  }h  i@  � s__n �@  :� s__c � 3  Z� m� \�a  �Y  ie:  `�� ���  ps:  z�  i�B  b�� ��  f�B  ]	�p�B  �� p�B  � p�B  @� kǞ
+   l"�  ��   �j�  pE�  �� p9�  �� p0�  �� l�:  ��   g`�  p;  �� p ;  �� p�:  �� v��   w;  ��   k��*�   q���D    yn  О   ���  ��  zh  i@  � {__n �@  �k�3�   Y�  ��  �  Zh  i@  V__c - 3  T\R'  /Y    e��  aN  �b   ���  X�  f��  � fȴ  �m� wմ  �� le:  ��   /n�  ps:  � jM:  ��   �p[:  � jt9  ��   -p�9  �    l�8  !�   2��  p�8  H� p�8  `�  lM:  &�   3͵  p[:  x� jt9  &�   -p�9  x�   i�;  (� 3M�  p�;  �� f�;  pt�v@�   p�;  �� f�;  pt���;  @�   �,�  f�;  pt� ��8  J�   �h�8  p�8  ��    k���    yt  `�d   �o�  ��  zh  i@  � {__c � 3  �g��  k�( �pȴ  �� p��  � m( wմ  W� le:  k�   /�  ps:  u� jM:  k�   �p[:  u� jt9  k�   -p�9  u�    l�8  ��   23�  p�8  �� p�8  ��  lM:  ��   3k�  p[:  �� jt9  ��   -p�9  ��   i�;  ��@ 3�  p�;  � p�;  :� v��   p�;  |� p�;  �� ��;  ��   �ʷ  p�;  ��  ��8  ��   �h�8  p�8  ��    k����     eFE  �   ПH   ��  �  pTE  �� p]E  �� phE  � ��A  ؟   �K�  p�A  0�  �.E  ߟX �ɸ  p<E  Z� l�;  �   ��  p�;  y�  j�;  �   �
<  f�;  p���8  �   d��8  f�8  p�   v�    phE  �� p]E  �� pTE  �� ����  ��0   ^�  � �  '�  Zh  i@  [�^  �'�   �7  e�  �l  �X   �G�  ��  f�  � f�  ��M:  #�p ���  f[:  �jt9  #�   -f�9  �  �FE  )�� �a�  hhE  p]E  �� pTE  �� ��A  )�   �ֹ  p�A  ��  �.E  3�� �6�  p<E  � j�;  p�   �
<  f�;  q���8  p�   d��8  f�8  q�   vP�   hhE  p]E  1� pTE  ^� k`���    ��@  ;�� �h�@  h�@  p�@  q�   ��  ��   ���   �  zh  i@  � u�^  < �  ��M:  ��� ��  p[:  �� gt9  ��� -p�9  ��   �M:  ��   �+�  p[:  �� jt9  ��   -p�9  ��   m� �__a �k   �oUY�  �M5  �FE  �� ��  hhE  p]E  �� pTE  ,� ��A  ��   䓻  p�A  ,�  �.E  ��0 ��  p<E  b� j�;   �   �
<  f�;  q���8   �   d��8  f�8  q�   v�    hhE  p]E  �� pTE  �� k���    �M:  ��   �<�  p[:  ��  �M:  ��   �Z�  p[:  ��  ��?  ��H ���  p�?    p�?  P  v��    p�?  n  p�?  �  ��?  ��` ���  p�?  �  p�?  �  �z8  ��` Vp�8  �  p�8  �  m` w�8  �     k۠z}    �E@  ��   �h\@  pS@  �     �7  eMG  ,Q  �   �@�  n�  f[G  � fdG  �����  �� � ���  r4*   �u   ��   !T   3   �E  �    �F  �  u\C  ��5  �u?)  ��  ��x �  �5# ��  ��e  �@  \R'  ��  ѽ  ��^  �Ľ  � ln;  2�
   �'�  px;   k8���   l�D  <�   �m�  pE  A j�@  <�   �h�@  p�@  m p�@  A   le:  B�   ���  ps:  �  ~x�   ��  pE  � lM:  x�   #��  p[:  �  j�?  }�   #p�?  � p�?  $ ���~  �Rug   kQ���  k^�eD  kg�3�   k���   �7  rn*  ��o   ���   !T   3   �E  �    �F  �  u\C  � 3  �u?)  ���  ��� ��  �5# ��  ��e  �@  ��^  �v�  � \R'  ���  ��  l�D  ��   ���  pE  7 j�@  ��   �h�@  p�@  c p�@  7   le:  ��   ��  ps:  �  ~�   ��  pE  � lM:  �   #J�  p[:  �  j�?  ��   #p�?  � p�?   ��~  �Rug   kǡ��  kء�D  k�3�   k��   �7  r�*  �L   ���   !T   3   �E  �    �F  �  u\C  P	��  �u?)  Q	��  ��� ��  ��^  S	�  � ~?�   z�  fE  ulM:  ?�   #D�  f[:  u j�?  D�   #p�?  ! p�?  N �S�~  �Ruw   �$�k/�3�   k\��   �7  �7  rp   `��   ��   ß  �,  ��|  |�,  a ��h  |�,  � �__a |�  ��H   �m� ��  �Y  � �__r ��7   �[F  v�� ���  pyF  q pnF  � ��E  v�� vp�E  q p�E  � �FB  v�� `pnB  � pbB  �    ��F  ��  �d�  p�F  " p�F  F p�F  � g�<  ��  �p�<  � p�<  � p�<  � g:  ��  �p@:   p4:  � p(:  � l�9  ��   iB�  p�9  X p�9  k p�9  ~ k���   j�8  â   gh�8  p�8  �     ��;  ��   ���  p�;    ��;  ��  ��  p�;  � p�;  � v�   f�;  Sf�;  W��;  �   ���  f�;  W ��8  �   �h�8  f�8  w s "#�   k��y    B6  oH  $ ��   �K�  fH  � f*H  �f5H  �f@H  ��8 h�  �JH  �UH  k�+   mP h@H  p5H   p*H  = pH  h mP wJH  � wUH  � ��G  #�p ���  p H  = p�G  h ��G  #�p vp�G  = p�G  h   ��<  3�� ���  p�<  M p�<  m p�<  � g:  3�� �p@:  � p4:  m p(:  � l�9  @�   i��  p�9  "	 p�9  5	 p�9  H	 kK��   j�8  c�   gh�8  p�8  [	    ��;  ;�   ���  p�;  �  ��;  N�� �?�  p�;  n	 p�;  �	 v��   f�;  Sf�;  W��;  ��   ��  f�;  W ��8  ��   �h�8  f�8  w s "#�   k3�y     ^�  � [�  ��  Zh  i@  [�^  ���  [%  �@  V__n �@   �7  eK�  �x ��T   ���  �  f[�  � fd�  �fp�  �f|�  ��t9  ��� ���  f�9  � ��:  ��   �A�  p;  �	 p ;  
 f�:  �v��   w;  G
 je:  ��   Ufs:  �   ��:  ��� �|�  f�:  r	�p�:  �
 f�:  �k��*   ��H  ��� ���  p�H   p�H  = p�H  P m� gpH  ��� �p�H   p�H  = p�H  P m� kǣH      ��@  ǣ   �h�@  p�@  s p�@  �   y�  �?   �-�  ��  zh  �9  �u%  �@  �{__n �@  �i�:   � ���  f�:  �	�p�:  � p�:  � le:   �   C��  ps:  �  k/��*   �� ^�  � ��  �  Zh  i@  [�^  ��  [%  �@  V__n �@  V__a ��   �7  B6  e��  �j 0�S   �'�  ��  f��  � f��  �f��  �f��  �f��  ��t9  5�  �m�  p�9    ��:  C�   ���  p;  % p ;  O p�:  � vC�   w;  � je:  C�   Ups:  �    ��:  S�8 ��  f�:  r	�p�:   f�:  �k���*   ��H  Y�   �~�  p�H  P p�H  d p�H  w vY�   jpH  Y�   �p�H  P p�H  d p�H  w vY�   kf�H      ��@  f�   �p�@  � p�@  � p�@  �   o�I   �  ���   ���  f�I  � f�I  �f�I  �f�I  ��P �  ��I  ��I  k��+   mh h�I  p�I  � p�I  � p�I    mh w�I  U w�I  � �]I  ä� ���  p{I  � ppI    �I  ä� vp-I  � p"I      �!=  Ӥ� �<�  pC=   p7=  % p+=  Z g:  Ӥ� �p@:  � p4:  % p(:  Z l�9  �   i�  p�9  � p�9  � p�9    k��   j�8  �   gh�8  p�8      ��;  ۤ   �Z�  p�;  �  ��;  �� ���  p�;  & p�;  g v �   f�;  Sf�;  W��;   �   ճ�  f�;  W ��8  )�   �h�8  f�8  w s "#�   kӤy     ^�  � ��  #�  Zh  i@  V__s ��5  V__n �@  V__a �#�   B6  e��  l 0�$   �C�  ��  f��  � f��  �f
�  �f�  ��.J  7�� ���  fYJ  �pMJ  � pAJ  � m� g�I  7�� �fJ  �p
J  � p�I  � m� kJ��I      ��@  J�   �f�@  �f�@  Pf�@  �   |(  �`��  ��  "�  zh  i@  � u%  �@  �t7i �@  � {__s ��5  �u<i �@  ��� �  �-  ��2   i�:  i�  ��  f�:  	�p�:  � p�:  M ie:  i�@ C��  ps:  � gM:  i�X �p[:  � gt9  i�X -p�9  �    kݦ�*   l�:  �   �I�  p;   p ;  m p�:  � v�   w;  Q   i�B  ��p ���  p�B  h p�B  � p�B  . p�B  x k̦
+   l�C  ��   ���  pD  � pD  H  �� D�  �Y�  ��%  �\iE  �� ���  pE  � iM:  �� #!�  p[:  � jt9  �   -p�9  �   j�?  �3   #p�?  � p�?  � v%�+   p�?   p�?  2 ��?  %�� ���  p�?  E p�?  Z �z8  %�� Vp�8  E p�8  Z m� w�8  o    kB�z}     lE  ߦ   �4�  fE  ud�lM:  ߦ   #��  f[:  ud� j�?  �   #p�?  � p�?  � ���~  �Ruc   ��k��C   �� �  Q  �@  � it9  c� �|�  p�9  !  i:  i�  ��  p@:  Y p4:  � p(:  � l�8  z�   g��  h�8  p�8  �  j�9  ��   ip�9  � p�9   p�9  ) k���    kc�*�   k���C   k���   y�   �"   �9�  ��  zh  i@  � u%  �@  �{__n �@  �u�^  ���  �le:  �   ���  fs:  �jM:  �   �f[:  �jt9  �   -f�9  �   k���   �7  y�  0�d   ���  �  }h  i@  < t�m �@  \ t7i �@  | t�^  ��  � t�m �@  � u<i �@  �i�:  7�@ ���  f;  �p ;  � p�:   m@ w;  = ge:  7�X Ups:   gM:  7�p �p[:   gt9  7�p -p�9        i�:  ]�� ��  f�:  	�p�:  � p�:  � k���*   q����   �7  y[  ��(   �1�  ��  zh  i@  � u%  �@  �u7i �@  �{__s ��5  �ln;  ��   ���  px;  � k����   kç��   elJ  V7  Ч   ���  Y�  fzJ  � p�J   f�J  �f�J  �f�J  �iFB  ԧ� +�  fnB  �!  fbB  �!   lFB  �   +2�  hnB  fbB  �!   ����  �� � ������  y�  �)   �p�  ��  zh  i@  � t��  �  . u�  �  �u�^  ��  �ie:  �� ��  ps:  M gM:  �� �p[:  M gt9  �� -p�9  M    jlJ  �   p�J  l p�J  � f�J  ��f�J  ��pzJ  � lFB  �   +h�  fnB  �K�  fbB  �A�   lFB  �   +��  hnB  fbB  �K�   k���    �7  y   �3   ���  ��  zh  i@  � t��  <�  � u�  <�  �{__s <�5  �ln;  /�	   ?�  fx;  �k8���   jlJ  8�   ?p�J   f�J  �f�J  ��f�J  ��fzJ  � lFB  <�   +�  fnB  �c�  fbB  �Y�   lFB  C�   +��  hnB  fbB  �c�   kL���    y~  `�%   ���  ��  zh  i@  � t��  v�    u�  v�  �u۶  vM5  �tnh  vM5  ? iFB  l�  {>�  fnB  ���  fbB  ��   lFB  z�   {d�  hnB  fbB  ���   �����  �� � ���  e�J  �9  ��%   ���  8�  f�J  � p�J  S f�J  �f�J  �pK  r iFB  �� ���  fnB  �"  fbB  �"   lFB  ��   ��  hnB  fbB  �"   �����  �� � ���  yJ  ��   �O�  D�  zh  i@  � t��  ��  � u�  ��  �{__l ��%  �g�J  Ĩ0 �fK  ��"�f�J  �p�J  � p�J  � f�J  � iFB  ĨH ���  fnB  �۰  fbB  �Ұ   lFB  Ҩ   ��  hnB  fbB  �۰   �ݨ��  �� � ������   y�  �%   �[�  �  zh  i@  � t��  ��  � u�  ��  �t۶  ��  � unh  ��  �iFB  �` ���  fnB  �  fbB  �   lFB  ��   ���  hnB  fbB  �   ����  �� � ���  y  �%   �-�  ��  zh  i@  � t��  ��   u�  ��  �t۶  ��  ; unh  ��  �iFB  �x ���  fnB  �\�  fbB  �l�   lFB  *�   ���  hnB  fbB  �\�   �5���  �� � ���  ^$  � ��  �  Zh  i@  V__s ��5  V__a ��   B6  e��  #o @�7   �:�  �  f��  � f�  �f�  ��n;  Q�   �y�  px;  Z kZ���   �.J  _�   ���  fYJ  �pMJ  m pAJ  � v_�   j�I  _�   �fJ  �p
J  m p�I  � v_�   kl��I      ��@  l�   �f�@  �f�@  Pf�@  �   ^�  � )�  K�  Zh  i@  V__l �%  V__a K�   B6  e�  �s ��$   �k�  ;�  f)�  � p2�  � f>�  ��.J  ��� ���  fYJ  �pMJ  � fAJ  �m� g�I  ��� �fJ  �p
J  � f�I  �m� k���I      ��J  ��   ��  f�J  �   ��@  ��   �f�@  �f�@  Pf�@  �   o�E  �t ��   �c�  f�E  � f�E  � rn2  ��   ���   {�  �5   �  �  u\C  /��  � u?)  0��  � K  K  Y�    ��  ��   f�  M5  Zh  i@  S�|  �M5  S�h  �M5  X__a ���   B6  e��  �i Щ    ��  ��   f�  M5  f��  � f��  �f��  �f��  ���H  ө   ��  f�H  �f�H  �f�H  �vө   jpH  ө   �f�H  �f�H  �f�H  �vө   k�H      ��@  �   �f�@  �f�@  Pf�@  �   Y�    ��  �   f�  �5  Zh  i@  S�|  �5  S�h  �5  X__a ��   B6  e��  �j �    �C�  ��   f�  �5  f��  � f��  �f�  �f�  ��.J  �   ���  fYJ  �fMJ  �fAJ  �v�   j�I  �   �fJ  �f
J  �f�I  �v�   k��I      ��@  �   �f�@  �f�@  Pf�@  �   Y�    �  A�   f�  �,  Zh  i@  S�|  �,  S�h  �,  X__a �A�   B6  e��  %h �    �j�  $�   f�  �,  f�  � f�  �f*�  �f5�  ���F  �   ���  f"G  �fG  ��f
G  ��v�   j�F  �   �f�F  �h�F  h�F  v�   k&���      ��@  &�   �f�@  �f�@  Pf�@  �   �U  =1�   [4  ��   >1�  �B  ?1�  ��  E]�   f4  �B   F]�  �C  G]�  �e  H]�  �8  I]�  ��  J]�  �

  X��   q4  ��  Y��  ��
  Z��  ��   `��  |4  ��  f��   �4  ��  g��  ��  h��  ��  n�   �4  ��	  o�  ��  p�  �H  vF�   �4  �`  wF�  �w  xF�  �   yF�  �~  �   �4  �   ��  ��  ��  �  ��  ��   ��  ��  ��  ��	  ��  ��  ���   �4  �  ���  �  ���  ��  ���  ��  ��   �4  ��  ��  ��  ��  ��  ��  �m  �Q�   �4  �	  �Q�  �2	  �Q�  ��  �Q�  �9  �Q�  �[  ���   �4  �J  ���  ��  ���  �7  ���  ��  ���   �4  �I	  ���  �$	  ���  ��   ���   �4  �N  ���  �p  ��   �4  ��  ��  �:  ��  ��  ��  �d   ��  ��  �a�    5  �  �a�  ��  �a�  ��	  э�   5  ��  ҍ�  �  ج�   5  ��  ٬�  ��  ڬ�  ��  ۬�  �+  ���   !5  ��  ���  ��   ���  �  ��   ,5  ��
  ��  ��  ��  �  �=�   75  �   �=�  �F  �=�  ��  �i�   B5  ��  �i�  ��  �i�  �D  O��   \5  ��  P��  �1  Q��  ��  W��   g5  �^  X��  ��  3��   r5  ��  4��  ��   8��   }5  ��  9��  �l	  =�  �5  �N  >�  �^  ?�  �L  @�  �a  DW�  �5  �B  EW�  ��	  FW�  �  GW�  �  HW�  �y  IW�  ��   ��   �5  ��  !��  ��*  �L  k �	�  #w �	�  �t �	�$  Zn �E��d  Z5   �  
Z5  
�5  
S5   ��O �O Z5  B�  
Z5  
�5  
�2   �us  s  Z5  d�  
Z5  
�2  
�2   ���  ��  �2  ��  
�5  
�5  
�2   �O2  Y2  �2  ��  
�5   ��`  �`  Z5  ��  
�5  
�2  
�2   5�  !��  Z5  ��  
W   	�  !�1  ��  
Z5   ��  Z5  �  
Z5   ��  �>  Y  
Z5    �Q   ��  ~ B{ �b �     �[ �x 
(0   �p  :   �  �x 
b%   (  _� �^   �  #  �� �  �  �   �  �  �   �  �O �   o  �O �   �	  pW   �   �  qW  !�   int   "�   �    #e   ` &�   ` '�   �^ (�   �^ )�   �T *�   �T +�   iY ,e   hY -�   �e 0�   �e 1�   [ 2�   [ 3�   Q 4�   Q 5�   �_ 6e   �_ 7�   �] :�   �] ;�   �Q >e   �Q ?�   s  Nx   �  Vx   .  <�   `  D�   �  W�   �  _�   �  e�   t   m�   a  u�     ~�   �  ��   3  ��   �  ��   H  ��   y  ��     ��   s  ��   T   ��   �  ��   F  ��   �  ��   �  ��     ��   V  ��   :   �  \	  2�   o  7�   �  <�   �  C�   �  �   	*  P  
�  �    rem �    +   +  	#@  �  
�  $L    rem %L    A  &[  std / �*  vP  w�  {�*  ��*  � +  �5+  �J+  ��+  ��+  ��+  ��+  ��+  �',  �G,  �h,  �s,  ��,  ��,  ��,  ��,  v  6�  x  K�  
�  M�   x  OT  _  �,  �   �  Qw  r  x  �,   �  R  �  �  �,     T8  �  �  �  �,   x  Z�  �  �,   x  \�  �  �,  -   x  _�  �  �,  �   x  c
    �,  	-   �  p�  -  -  8  �,  -   �  t�  -  P  [  �,  	-   �  {k  v  �,  �    n	 ~%  �  �  �,  -   �  ��  -  �  �  �,   �  �h  -  �  �,    -   :-  �  �s   � �  �S L%  &0@i1  �=  ��  �b  �:   Fe  ��   �3  �=  B  t1  z1      eq �<-  -  d  z1  z1    lt ��1  -  �  z1  z1   !��  eF  �   �  �1  �1  �   !�K  �9  �  �  �1   !�(  
!  �1  �  �1  �  z1   !1  �A  �1    �1  �1  �   !�5  �'  �1  +  �1  �1  �   !�3  �A  �1  O  �1  �     !+  :    i  �1     !�C   �P    �  z1   !�B  $6  -  �  �1  �1   "eof (�:    #?  ,N0    �1    _� �^   0�   1�   2�   3�   5Y  6o  7�  8�  :  ;  <-  =C  ?�  @�  Bx   C�   D�   E�   Gd  Hz  I�  J�  L  M"  N8  ON  Q�  R�  G�  c�?  �L   K  \0	  $B-   %�e  _�  %�4  c�1  %�J  d�1  ��  q�  �  �1   ��  s	  	  �1  �1   &W  y$	  �1  �     �  5�1  6�2  73  �J  pr"  '�B  �	  (�   )%  �   *�B  �	  �	  23  �  �1   +�B  �	  23  �     %�e  y�  ,[V  �	  �	  )�G  !V	   %<  x�  %�4  {�  %�J  |�  %�J  �.  %`S  ��0  %~J  �}"  %�J  ��"  �%  �[
  
�K  ��	   
I  ��	  
:!  �"3   %H  �  (*
   -�3  2�	  -�G  7+  -t3  Bb3  .�'  ��O  J3  V  ��N  -  �
  �
  m3   3  �o+  -  �
  �
  m3   �P  ��O  �
  �
  D3   �M  ��P    	  D3   �,  �-    '  D3  �	   �+  ��R  �  >  D  D3   3  �   �  [  k  D3  �1  �1   !�/  !�B  D3  �  �	  �	  �1   �O  �|6  �  �  D3  �1   /(  ��6  �  �  D3  �1   0�   �-  �  �  �  D3   1�1  o�*  �  �  D3  �1  �	    0�A  $n%  �  '  -  83   0�A  (�I  �  E  P  >3  �   0"A  ,�%  D3  h  n  83   0�1  2E)  �	  �  �  83   0�/  6;&  �	  �  �  83   /�>  :�>  �  �  >3   0S  A:2  �	  �  �  83  �	  +   /�#  K�(       83  �	  �	  +   09  S>$  �	  -  =  83  �	  �	   0-U  [�7  -  U  `  83  +   2�5  d�-  �  �  +  �	   2	1  m�P  �  �  +  �	   2�3  v\-  �  �  �	  :    2nU  ��-  �  �  �	  �	   2nU  �nG     �  
  
   2nU  ��      �  �  �   2nU  �IP  @  �  +  +   !�J  �rR  �   _  �	  �	   /�=  ��H  s  �  >3  �	  �	  �	   /V  �)  �  �  >3   3�'  �D*  J3  4�0  ��  �  >3   5�0  ��  �  >3  �1   4�0  ��    >3  P3   4�0  �  '  >3  P3  �	  �	   4�0  �8  R  >3  P3  �	  �	  �1   4�0  �c  x  >3  +  �	  �1   4�0  ��  �  >3  +  �1   4�0  ��  �  >3  �	  :   �1   4�0   �  �  >3  V3   4�0  �  �  >3  �"  �1   4�0  "    >3  �    6�  *,Q  \3  1  <  >3  P3   6�  2�G  \3  U  `  >3  +   6�  =�%  \3  y  �  >3  :    6�  Mo_ \3  �  �  >3  V3   6�  Y.c \3  �  �  >3  �"   6S� f�&  �	  �  �  >3   6S� q�>  
    
  83   7end y<  �	  #  )  >3   7end �6;  
  B  H  83   6I ��$  
  a  g  >3   6I ��7  
  �  �  83   6��  �lC  
  �  �  >3   6��  �CM  
  �  �  83   6)^ �^\ 
  �  �  83   6%] ��a 
  �    83   6hf �*] 
    !  83   6wY �Je 
  :  @  83   6r ��R  �	  Y  _  83   6�K  �r5  �	  x  ~  83   6�3  �j=  �	  �  �  83   8�� ��  �  �  >3  �	  :    8�� ��F  �  �  >3  �	   8be  VT �  �  >3   6I  v  �	      83   8�E  &|U  1  <  >3  �	   8�1  -�  Q  W  >3   6�� 5�?  -  p  v  83   6�:  D�6  �	  �  �  83  �	   6�:  UW  �	  �  �  >3  �	   7at k
/  �	  �  �  83  �	   7at ��7  �	  �    >3  �	   6��  ��O �	    #  >3   6��  �}Y �	  <  B  83   6�G  �@\ �	  [  a  >3   6�G  �e �	  z  �  83   6�F  ��/  \3  �  �  >3  P3   6�F  �k:  \3  �  �  >3  +   6�F  ��H  \3  �  �  >3  :    6�F  �x` \3      >3  �"   6@  �A:  \3  )  4  >3  P3   6@  ��1  \3  M  b  >3  P3  �	  �	   6@  ��D  \3  {  �  >3  +  �	   6@  ��*  \3  �  �  >3  +   6@  �6  \3  �  �  >3  �	  :    6@  �] \3  �  �  >3  �"   8�G  -aN      >3  :    6�3  <b*  \3  5  @  >3  P3   6�3  Ipf \3  Y  d  >3  V3   6�3  ^ 2  \3  }  �  >3  P3  �	  �	   6�3  n�=  \3  �  �  >3  +  �	   6�3  z�T  \3  �  �  >3  +   6�3  � @  \3  �    >3  �	  :    6�3  ��a \3  !  ,  >3  �"   8� ��E  A  V  >3  �	  �	  :    8� ��V k  {  >3  �	  �"   6� �\+  \3  �  �  >3  �	  P3   6� �u>  \3  �  �  >3  �	  P3  �	  �	   6� |=  \3  �    >3  �	  +  �	   6� "�@  \3    .  >3  �	  +   6� 9k<  \3  G  \  >3  �	  �	  :    6� K�'  �	  u  �  >3  �	  :    6bL  d�R  \3  �  �  >3  �	  �	   6bL  t�2  �	  �  �  >3  �	   6bL  �L&  �	  �  �  >3  �	  �	   8H�  �M\     >3   6�%  �9F  \3  /  D  >3  �	  �	  P3   6�%  �|<  \3  ]  |  >3  �	  �	  P3  �	  �	   6�%  ��T  \3  �  �  >3  �	  �	  +  �	   6�%  ��A  \3  �  �  >3  �	  �	  +   6�%  b>  \3  �    >3  �	  �	  �	  :    6�%  3%  \3  )  >  >3  �	  �	  P3   6�%  'V7  \3  W  q  >3  �	  �	  +  �	   6�%  <�+  \3  �  �  >3  �	  �	  +   6�%  Q'S  \3  �  �  >3  �	  �	  �	  :    6�%  vj.  \3  �    >3  �	  �	  �  �   6�%  ��9  \3    8  >3  �	  �	  +  +   6�%  �C  \3  Q  k  >3  �	  �	  �	  �	   6�%  �>/  \3  �  �  >3  �	  �	  
  
   6�%  �b \3  �  �  >3  �	  �	  �"   0�?  ��&  \3  �  �  >3  �	  �	  �	  :    0�1  �O  \3    0  >3  �	  �	  +  �	   !,)  �z-  �  T  �	  :   �1   !+E  �3J  �  x  �	  :   �1   6�5  �)  �	  �  �  83  �  �	  �	   8n	 @D  �  �  >3  \3   6W�  �6  +  �  �  83   6�A  %�A  +  �    83   6��  ,Z5  �	    #  83   6�(  <;  �	  <  Q  83  +  �	  �	   6�(  I�%  �	  j  z  83  P3  �	   6�(  X�5  �	  �  �  83  +  �	   6�(  i^   �	  �  �  83  :   �	   6�(  v�S  �	  �  �  83  P3  �	   6�(  �K  �	    #  83  +  �	  �	   6�(  �o?  �	  <  L  83  +  �	   6�(  �J5  �	  e  u  83  :   �	   6NW  ��Q  �	  �  �  83  P3  �	   6NW  ��I  �	  �  �  83  +  �	  �	   6NW  ��,  �	  �  �  83  +  �	   6NW  ��;  �	      83  :   �	   6�S  ��I  �	  7  G  83  P3  �	   6�S  T?  �	  `  u  83  +  �	  �	   6�S  05  �	  �  �  83  +  �	   6�S  $S:  �	  �  �  83  :   �	   6�>  2hL  �	  �  �  83  P3  �	   6�>  CUB  �	  	      83  +  �	  �	   6�>  Q�2  �	  7   G   83  +  �	   6�>  b�K  �	  `   p   83  :   �	   6�4  qT  �	  �   �   83  P3  �	   6�4  ��K  �	  �   �   83  +  �	  �	   6�4  ��5  �	  �   �   83  +  �	   6�4  �N.  �	  	!  !  83  :   �	   6U+  �)  J	  2!  B!  83  �	  �	   6��  �!1  �   [!  f!  83  P3   6��  ��T  �   !  �!  83  �	  �	  P3   6��  ��O  �   �!  �!  83  �	  �	  P3  �	  �	   6��  	;.  �   �!  �!  83  +   6��  (	�B  �   	"  "  83  �	  �	  +   6��  C	�,  �   7"  Q"  83  �	  �	  +  �	   [
  9!T  :   :�E    :�F  �   � >J	  �&  �7  J	  Qf /l#  %�J  6+  
t :�"   %�e  5�  
�x ;�"  %`S  7+  ;�w >�"  �"  �3  �"  �"   �w B#  	#  �3   r G�i �"  !#  '#  �3   S� K�m �"  ?#  E#  �3   <end O;u �"  ]#  c#  �3   =_E :    q#  Y� �x w�$  >~ ��    >z �s3  ;�x y�#  �#  y3   ;�x |�#  �#  y3  �   3   �3  �Nz �#  �#  y3  �   3   �1  ��y $  $  y3   ~ ��� �   #$  )$  �3   �| ��| 3  @$  F$  �3   } ��y �$  ]$  c$  �3   9� ��y r"  z$  �$  �3   ?�  �� -  �$  �3    v#  �� Ĭ%  
~ ��    
z �s3  �� ��$  �$  �3   �� ��$  �$  �3  �   3   �3  ҁ{ %  %  �3  �   3   �1  ��} 1%  7%  �3   ~ ��{ �   O%  U%  �3   �| �} 3  m%  s%  �3   9� ��x r"  �%  �%  �3   @�  �y -  �%  �3    �"  �$  � 'A��  )�   <�3   =�3   >�3   @I4   AT4   Bn4   C�4   D�4   E�4   F�4   G�4   H5  Gz !<<&  B_V2 !�C!�+&   Ayy "aAo� "dA� "h#P�0  #Q�0  #R�0  #S�0  #T�0  D�~ @�&  E�| E�y E�~ E  Q� $)�'  F�~ $1'  E }  E�} E�} E�� Ej| E�| E[| E�} Ey| EDy 	E{ 
E_ ESy  G} $C'   �&  G�} $F'  G�} $L'  G�� $O'  Gm| $R'  G�| $U'  G^| $X'  G�} $['  G|| $a'  GGy $g'  	G{ $l'  
Gb $r'  GVy $x'   ד  %��'  ��  %��  � %��  �4  %��1  9{�  �   H�� �'  &�� ?�'  6    H�z (  &�z L(  �6    Hz 2(  &z 9+(  �6    H��  N(  &��  �G(  �6    Hv� j(  &v� �c(  �6    H� �(  I� }(  "7    J�x Rv#  �(  z&   K�z 6�~ Kz :-| K	@  >�N  K�} BG} �p F]u �(  +   � J)} �(  +   }� N� )  +   � R� )  +   }z VA .)  +   ��  Z)�  D)  +  L �8 j#< Y)  +    ns n)  +   by r"{ �)  +   �{ v�z �)  +   t4 z�/ �)  +   H| �)  M| >�)  ?G  v#    | ~�| �)  �    HN| *  NN| c�)  �H  v#    F| �� *  �    K � �a} | ��z :*  �&   O	[ OG*   �  P%�  e �  [*  �  O6y )m*   �%  QIc  1�*   �%  Q& "j�*   <&  Q�~ "k�*   E&  Q{ "l�*   N&  .�| ny 3  .1 N�{ 3   J� ��   �*  �*   �*  RJ�  >+  +  +   �� +  :   J�  H�   5+  +   J�  IL   J+  +   J�  ��  s+  s+  s+  S   S   z+   y+  S�+  T�   �+  s+  s+   Udiv P  �+  �   �    J    ��  �+  +   V�   �  �+  L   L    V�  .�   �+  +  S    V�  \S   ,  ,  +  S     ,    V3  >�   G,  ,  +  S    W�  h,  �  S   S   z+   Xk� q�   Y�  |�,  �    J  W+  �,  +  �,   �  J  fL   �,  +  �,  �    J�  g^   �,  +  �,  �    J?  ��   �,  +   -  �  Z�  [-  Z-  �  �  $   �G1  �  '$(,�  (-�  K  (:�.  %�e  (=�  %� (?�  %"  (@+  %�4  (A�1  %�J  (B�1  �A  (O�-  �-  �1   �A  (Q�-  �-  �1  �1   �A  (V�-  �-  �1  �    �
 (Y51  Z-  �-  �-  �1  r-   �
 (]�R  f-  .  .  �1  ~-   � (c?  Z-  4.  D.  �1  N-  s+   _ (m.   X.  h.  �1  Z-  N-   �3  (q89  N-  �.  �.  �1   =_Tp :    B-  \ZD  )��0  ]F�  )��   ^��  )��'  ^�4  )��'  ^� )��'  4��  )��.  �.  25   5��  )��.  
/  25  85   6*  )��}  �.  #/  )/  C5   6Ư  )�?s  �.  B/  H/  C5   6�F  )�Ϭ  I5  a/  g/  25   6�F  )��  �.  �/  �/  25  �    6a�  )�
�  I5  �/  �/  25   6a�  ) ��  �.  �/  �/  25  �    6�:  ),�  �.  �/  �/  C5  �.   6�F  )		n  I5  0  0  25  �.   6(*  )��  �.  /0  :0  C5  �.   6 I  )h�  I5  S0  ^0  25  �.   6�O  )7k  �.  w0  �0  C5  �.   6WC  )]�  85  �0  �0  C5   9{�  �  9�  J	   8E  F*; *1�0  E�8  E�; EN;  G�= *5�0   �0  �.  _U  A"3  1  O5  �    _9+  N"3  "1  O5  �    `A� -z �   �  �  +  A     �� 2*  &7a1  a&8�   b+pO qO +!a1  Z  ZB  B    Zi  Ye �[ Z:   Z+  B-  Z�.  �.  �  Z0	  �  8,�2  
�{  ,�   
]�  ,�  
\�  , �  
�D  ,!�  
�3  ,"�  
U>  ,#�  
&�  ,$�  
�  ,%�  
�*  ,&�   
ڡ  ,':   $
�U  ,(:   %
TL  ,):   &
�I  ,*:   '
Q  ,+:   (
�C  ,,:   )
�J  ,-:   *
1  ,.�  ,
o(  ,/:   0
�U  ,0:   1
PL  ,1:   2
�I  ,2:   3
Q  ,3:   4
�C  ,4:   5
�J  ,5:   6 J)%  ,K�  3  �   +   XGT  ,P3  �1  �  - �   �   V	  �"  J	  [
  Z[
  Z�"  [J	  ZJ	  c^   m3  d Q"  l#  v#  Zl#  �$  �"  �%  �$  �%  �l  .L   j�  .#L   etm ,.,I4  
,g  ..�    
�  ./�   
�  .0�   
��  .1�   
��  .2�   
��  .3�   
��  .4�   
�  .5�   
d�  .6�    
��  .7L   $
~�  .8+  ( X\�  .>�3  Jѯ  .H+  n4  �3  �3   J��  .M�3  �4  �4   �3  J�  .C�3  �4  �4   �3  J#�  .a�  �4  �4   �4  �3  J�� .f�  �4  �4   �4  �3  J��  .W�4  �4  �4   J[v  .\�4  5  �4   J��  .RS   25  �  S   +  �4   �.  Z>5  �  �0  Z�.  "3  f�0  �5  gXF  AO5  g\;  A�   hi�T  C"3    j  �5  �5  kh  �5   83  f�
  �5  hl__p ��    f1  �5  gXF  NO5  g\;  N�    j�  �5  �5  kh  �5  m__a �6   D3  �1  �'  j�'  6  $6  kh  $6   6  j$  76  A6  kh  A6   �3  j)$  T6  ^6  kh  A6   j�#  l6  �6  kh  �6  m__v |�   g=8 |�6   y3  3  �'  j(  �6  �6  kh  �6   �6  (  j(  �6  �6  kh  �6   �6  2(  j;(  �6  �6  kh  �6   �6  N(  jW(  7  7  kh  7   �6  j(  ns(  	�97  C7  kh  C7   "7  j�-  V7  `7  kh  `7   �1  j�  s7  }7  kh  }7   �1  j�-  �7  �7  kh  `7  k#  -3   j	  �7  �7  kh  }7  k#  -3   j�-  �7  �7  kh  `7  �7   �1  j�  �7  	8  kh  }7  m__a s	8   �1  j  8  &8  kh  �5   jP  48  >8  kh  �5   n�	  O8  b8  kh  b8  k#  -3   23  j�  u8  �8  kh  �8  k#  -3   >3  jc$  �8  �8  kh  A6   f�(  �8  g2� Rz&   o�5  0�$   ��8  ?9  p�5  � p�5  5 q�5  4�8 �59  r�5  p�5  o sU5  4�8 Vrj5  p_5  o t8 uv5  �    vO��   w�(  `�#   ��9  x�6  m�   7o9  p�6  �  vj�=Q  v��QQ   w�(  ��#   ��9  x�6  ��   ;�9  p�6  �  v��=Q  v��QQ   w�(  ��#   �:  x�6  ͪ   ?�9  p�6     vʪ=Q  v�QQ   w�(  �#   �K:  x7  ��   C8:  p7  "   v��=Q  v�QQ   w�(   ��   �z;  y__s F+  � qg8  M�P G�:  pu8  5  z&8  M�p #�:  p48  5   {�5  V�� #p�5  H  p�5  ]  |x��8  }Rus   xg8  ��   GI;  ~u8  ut�&8  ��   #;  ~48  ut� ��5  ��   #p�5  {  p�5  �  |���8  }Rus   v2�=Q  �D��M�vp�QQ  v��}Q  v���Q   w�(  ���   ��<  y__s J+  � qg8  ݫ� K	<  pu8  �  z&8  ݫ� #�;  p48  �   {�5  �� #p�5  �  p�5  �  |��8  }Rus   xg8  �   Kx<  ~u8  ut�&8  �   #C<  ~48  ut� ��5  %�   #p�5  ! p�5  .! |4��8  }Rus   v«=Q  �ԫ�ݫv �QQ  v�}Q  v��Q   w�(  @��   ��=  y__s N+  � qg8  m�� O8=  pu8  A! z&8  m� #=  p48  A!  {�5  v�( #p�5  T! p�5  i! |���8  }Rus   xg8  ��   O�=  ~u8  ut�&8  ��   #r=  ~48  ut� ��5  ��   #p�5  �! p�5  �! |Ĭ�8  }Rus   vR�=Q  �d��m�v��QQ  v��}Q  v���Q   w)  Ь�   �?  y__s R+  � qg8  ��@ Sg>  pu8  �! z&8  ��` #3>  p48  �!  {�5  �x #p�5  �! p�5  �! |(��8  }Rus   xg8  ?�   S�>  ~u8  ut�&8  ?�   #�>  ~48  ut� ��5  E�   #p�5  " p�5  :" |T��8  }Rus   v�=Q  ������v �QQ  v5�}Q  v=��Q   w)  `��   �6@  y__s V+  � qg8  ��� W�?  pu8  M" z&8  ��� #b?  p48  M"  {�5  ��� #p�5  `" p�5  u" |���8  }Rus   xg8  ϭ   W@  ~u8  ut�&8  ϭ   #�?  ~48  ut� ��5  խ   #p�5  �" p�5  �" |��8  }Rus   vr�=Q  ������v��QQ  vŭ}Q  vͭ�Q   w.)  ��   ��A  �-  Z+  � L����   �A  iR'  \�%  �a� _�%  �" �__s `>5  �" ��| aA   �# qg8  O�� eA  pu8  $ z&8  O�  #�@  p48  $  {�5  X� #p�5  $ p�5  A$ |z��8  }R�k   xg8  ��   eA  ~u8  �l�&8  ��   #JA  ~48  �l� ��5  ��   #p�5  _$ p�5  �$ |���8  }R�k   v��Q  v'�"1  v3�=Q  �F��O�vr�QQ  v��}Q   v���Q   wD)  ���   ��B  y__s j+  � qg8  ݮ0 kRB  pu8  �$ z&8  ݮP #B  p48  �$  {�5  �h #p�5  �$ p�5  �$ |��8  }Rus   xg8  �   k�B  ~u8  ut�&8  �   #�B  ~48  ut� ��5  %�   #p�5  �$ p�5  % |4��8  }Rus   v®=Q  �Ԯ�ݮv �QQ  v�}Q  v��Q   wY)  @��   �!D  y__s n+  � qg8  m�� o�C  pu8  %% z&8  m�� #MC  p48  %%  {�5  v�� #p�5  8% p�5  M% |���8  }Rus   xg8  ��   o�C  ~u8  ut�&8  ��   #�C  ~48  ut� ��5  ��   #p�5  k% p�5  �% |į�8  }Rus   vR�=Q  �d��m�v��QQ  v��}Q  v���Q   wn)  Я�   �PE  y__s r+  � qg8  ��� s�D  pu8  �% z&8  ��� #|D  p48  �%  {�5  � #p�5  �% p�5  �% |(��8  }Rus   xg8  ?�   sE  ~u8  ut�&8  ?�   #�D  ~48  ut� ��5  E�   #p�5  �% p�5  & |T��8  }Rus   v�=Q  ������v �QQ  v5�}Q  v=��Q   w�)  `��   �F  y__s v+  � qg8  ��  w�E  pu8  1& z&8  ��@ #�E  p48  1&  {�5  ��X #p�5  D& p�5  Y& |���8  }Rus   xg8  ϰ   wNF  ~u8  ut�&8  ϰ   #F  ~48  ut� ��5  հ   #p�5  w& p�5  �& |��8  }Rus   vr�=Q  ������v��QQ  vŰ}Q  vͰ�Q   w�)  �m   �?G  y__s z+  � qg8  �p {G  pu8  �& z&8  �� #�F  p48  �&  {�5   �� #p�5  �& p�5  �& |H��8  }Rus   v�=Q  ����v@�QQ  vU�}Q  v]��Q   �)  j�)  SG  jG  kh  jG  ��} >v#   ?G  ��)  `��   ��H  y__i ~�   � qEG  |�� ��H  p\G  �& ~SG  S�8  |�   ?�G  ~�8  ��	   zg8  ��� ?DH  pu8  S' z&8  �� #H  p48  S'  {�5  ��( #p�5  h' p�5  }' |ͱ�8  }Ruc   g8  �   ?�H  ~u8  ud�&8  �   #H  ~48  ud� ��5  �   #p�5  �' p�5  �' |���8  }Ruc   ��� vs�=Q  vz��*  vűQQ  vڱ}Q  v��Q   �)  j�)  �H  I  kh  I  g�} cv#   �H  w*   ��   ��J  y__i ��   � q�H  �@ �EJ  pI  �' ~�H  Sqg8  7�x d�I  pu8  ( z&8  7�� #�I  p48  (  {�5  @�� #p�5  ( p�5  -( |q��8  }Rub   xg8  ��   d8J  ~u8  ud�&8  ��   #J  ~48  ud� ��5  ��   #p�5  K( p�5  x( |���8  }Rub   �.��7� x�8  �   �jJ  ~�8  uv��*   v�=Q  vi�QQ  v~�}Q  v���Q   w*  ��#   ��J  x(7  ��   ��J  p97  �(  v��=Q  vòQQ   w%*  вB   �K  �~ ��&  � v߲=Q  ��v��QQ  v
�}Q  v��Q   �D  O,K   �  ��  P,K  �1  Q,K  ��  WXK   �  �^  XXK  �U  =wK   �  ��   >wK  �B  ?wK  ��  E�K      �B   F�K  �C  G�K  �e  H�K  �8  I�K  ��  J�K  �

  X�K     ��  Y�K  ��
  Z�K  ��   `"L    ��  f4L   !  ��  g4L  ��  h4L  ��  n`L   ,  ��	  o`L  ��  p`L  �H  v�L   7  �`  w�L  �w  x�L  �   y�L  �~  �L   B  �   ��L  ��  ��L  �  ��L  ��   ��L  ��  ��L  ��	  ��L  ��  �%M   M  �  �%M  �  �%M  ��  �%M  ��  �^M   X  ��  �^M  ��  �^M  ��  �^M  �m  ��M   c  �	  ��M  �2	  ��M  ��  ��M  �9  ��M  �[  ��M   n  �J  ��M  ��  ��M  �7  ��M  ��  �N   y  �I	  �N  �$	  �N  ��   �BN   �  �N  �BN  �p  �aN   �  ��  �aN  �:  �aN  ��  �aN  �d   �aN  ��  ɧN   �  �  ʧN  ��  ˧N  ��	  ��N   �  ��  ��N  �  ��N   �  ��  ��N  ��  ��N  ��  ��N  �+  �+O   �  ��  �+O  ��   �+O  �  �WO   �  ��
  �WO  ��  �WO  �  �O   �  �   �O  �F  ��O  ��  �O   �  ��  ��O  ��  ��O  ��  3�O   �  ��  4�O  ��   8�O   �  ��  9�O  �l	  =P  
  �N  >P  �^  ?P  �L  @P  �a  DRP    �B  ERP  ��	  FRP  �  GRP  �  HRP  �y  IRP  ��   �P      ��  !�P  ��0   �:*  �`*  �r*  ��*  ��*  ��*  �'   �'  �"'  �.'  �:'  �F'  �R'  �^'  �j'  �v'  	��'  
��'  ��'  ��  �  QQ  ^    ��  kQ  �  �  kQ   qQ  �}Q  �   �  �Q  �   �>  Y  �Q  �   �O2  Y2  ^   +    �1   <�  1� �� �b �     �e std  H   v  6�  x  K�  �  MH    x  Ob   m   J   H    	�  Qw  �   �   J    	�  R  �   �   J    
  T8  H   �   �   P    x  Z�   �   J    x  \�   �   J   V    x  _�     J   �   x  c  #  J   a    �  p�  g   ;  F  J   V    �  t�  g   ^  i  J   a    �  {y  �  J   m    n	 ~%  �  �  J   g    �  ��  t   �  �  P    �  �h  {   �  P     ;    :;   �  �\   � �  �S L%  0@7%  �=  ��  �b  �"  Fe  �m   �3  �=  P  B%  H%      eq �<-  t   r  H%  H%   lt ��1  t   �  H%  H%   ��  eF  m   �  N%  N%  �   �K  �9  �  �  N%   �(  
!  N%  �  N%  �  H%   1  �A  T%    T%  N%  �   �5  �'  T%  9  T%  N%  �   �3  �A  T%  ]  T%  �      +  :     w  Z%   +  �C   �P  +  �  H%   �B  $6  t   �  Z%  Z%   eof (�:  +  ?  ,N0  +  Z%    _� �D"  0�"  1�"  2�"  3�"  5M#  6c#  7y#  8�#  :�"  ;#  <!#  =7#  ?�#  @�#  B�"  C�"  D�"  E�"  GX#  Hn#  I�#  J�#  L #  M#  N,#  OB#  Q�#  R�#  �?  �`"  K  	\6  �    �e  	_�  �4  	cn%  �J  	dt%  ��  	q�    �%   ��  	s    �%  �%   W  	y*  �%  m     �  
5�%  
6�&  
7�&  �J  px  �B  �   �   !%  �$   "�B  �  �  '  �$  �%   #�B  �  '  m     �e  y�  $[V  �  �  !�G  !\   <  x�  �4  {�  �J  |�  �J  �!  `S  ��!  ~J  �x  �J  �}  �%  �a  �K  ��   I  ��  :!  ��&   %H  �   0   %�3  2�  %�G  7*%  %t3  B7'  &�'  ��O  '  
V  ��N  t   �  �  B'   
3  �o+  t   �  �  B'   	�P  ��O  �  �  '   	�M  ��P  	    '   	�,  �-  "  -  '  �   
�+  ��R  �$  D  J  '   
3  �   �$  a  q  '  �%  �%   �/  !�B  '  �  �  �  �%   	�O  �|6  �  �  '  �%   '(  ��6  �  �  '  �%   (�   �-  �$  �  �  '   )�1  o�*  �$    '  �%  �    (�A  $n%  �$  -  3  '   (�A  (�I  �$  K  V  '  �$   ("A  ,�%  '  n  t  '   (�1  2E)     �  �  '   (�/  6;&     �  �  '   '�>  :�>  �  �  '   (S  A:2  �  �  �  '  �  $%   '�#  K�(  	  	  '  �  �  $%   (9  S>$  �  3	  C	  '  �  �   (-U  [�7  t   [	  f	  '  $%   *�5  d�-  �	  �$  $%  �   *	1  m�P  �	  �$  $%  �   *�3  v\-  �	  �$  �  �"   *nU  ��-  �	  �$         *nU  �nG  
  �$       *nU  ��   &
  �$  �$  �$   *nU  �IP  F
  �$  $%  $%   �J  �rR  m   e
  �  �   '�=  ��H  y
  �
  '  �  �  �   'V  �)  �
  �
  '   +�'  �D*  '  ,�0  ��
  �
  '   -�0  ��
  �
  '  �%   ,�0  ��
    '  %'   ,�0  �  -  '  %'  �  �   ,�0  �>  X  '  %'  �  �  �%   ,�0  �i  ~  '  $%  �  �%   ,�0  ��  �  '  $%  �%   ,�0  ��  �  '  �  �"  �%   ,�0   �  �  '  +'   ,�0  �    '  �  �%   ,�0  "    '  m    .�  *,Q  1'  7  B  '  %'   .�  2�G  1'  [  f  '  $%   .�  =�%  1'    �  '  �"   .�  Mo_ 1'  �  �  '  +'   .�  Y.c 1'  �  �  '  �   .S� f�&     �  �  '   .S� q�>    
    '   /end y<     )  /  '   /end �6;    H  N  '   .I ��$  $  g  m  '   .I ��7    �  �  '   .��  �lC  $  �  �  '   .��  �CM    �  �  '   .)^ �^\   �  �  '   .%] ��a       '   .hf �*]   !  '  '   .wY �Je   @  F  '   .r ��R  �  _  e  '   .�K  �r5  �  ~  �  '   .�3  �j=  �  �  �  '   0�� ��  �  �  '  �  �"   0�� ��F  �  �  '  �   0be  VT �    '   .I  v  �    "  '   0�E  &|U  7  B  '  �   0�1  -�  W  ]  '   .�� 5�?  t   v  |  '   .�:  D�6  �  �  �  '  �   .�:  UW  �  �  �  '  �   /at k
/  �  �  �  '  �   /at ��7  �  �  
  '  �   .��  ��O �  #  )  '   .��  �}Y �  B  H  '   .�G  �@\ �  a  g  '   .�G  �e �  �  �  '   .�F  ��/  1'  �  �  '  %'   .�F  �k:  1'  �  �  '  $%   .�F  ��H  1'  �  �  '  �"   .�F  �x` 1'      '  �   .@  �A:  1'  /  :  '  %'   .@  ��1  1'  S  h  '  %'  �  �   .@  ��D  1'  �  �  '  $%  �   .@  ��*  1'  �  �  '  $%   .@  �6  1'  �  �  '  �  �"   .@  �] 1'  �    '  �   0�G  -aN    "  '  �"   .�3  <b*  1'  ;  F  '  %'   .�3  Ipf 1'  _  j  '  +'   .�3  ^ 2  1'  �  �  '  %'  �  �   .�3  n�=  1'  �  �  '  $%  �   .�3  z�T  1'  �  �  '  $%   .�3  � @  1'  �    '  �  �"   .�3  ��a 1'  '  2  '  �   0� ��E  G  \  '     �  �"   0� ��V q  �  '     �   .� �\+  1'  �  �  '  �  %'   .� �u>  1'  �  �  '  �  %'  �  �   .� |=  1'  �    '  �  $%  �   .� "�@  1'  $  4  '  �  $%   .� 9k<  1'  M  b  '  �  �  �"   .� K�'     {  �  '     �"   .bL  d�R  1'  �  �  '  �  �   .bL  t�2     �  �  '      .bL  �L&     �    '         0H�  �M\     '   .�%  �9F  1'  5  J  '  �  �  %'   .�%  �|<  1'  c  �  '  �  �  %'  �  �   .�%  ��T  1'  �  �  '  �  �  $%  �   .�%  ��A  1'  �  �  '  �  �  $%   .�%  b>  1'  �    '  �  �  �  �"   .�%  3%  1'  /  D  '        %'   .�%  'V7  1'  ]  w  '        $%  �   .�%  <�+  1'  �  �  '        $%   .�%  Q'S  1'  �  �  '        �  �"   .�%  vj.  1'  �    '        �$  �$   .�%  ��9  1'  $  >  '        $%  $%   .�%  �C  1'  W  q  '               .�%  �>/  1'  �  �  '             .�%  �b 1'  �  �  '        �   (�?  ��&  1'  �    '  �  �  �  �"   (�1  �O  1'    6  '  �  �  $%  �   ,)  �z-  �$  Z  �  �"  �%   +E  �3J  �$  ~  �  �"  �%   .�5  �)  �  �  �  '  �$  �  �   0n	 @D  �  �  '  1'   .W�  �6  $%  �  �  '   .�A  %�A  $%    
  '   .��  ,Z5  �  #  )  '   .�(  <;  �  B  W  '  $%  �  �   .�(  I�%  �  p  �  '  %'  �   .�(  X�5  �  �  �  '  $%  �   .�(  i^   �  �  �  '  �"  �   .�(  v�S  �  �  �  '  %'  �   .�(  �K  �    )  '  $%  �  �   .�(  �o?  �  B  R  '  $%  �   .�(  �J5  �  k  {  '  �"  �   .NW  ��Q  �  �  �  '  %'  �   .NW  ��I  �  �  �  '  $%  �  �   .NW  ��,  �  �  �  '  $%  �   .NW  ��;  �    $  '  �"  �   .�S  ��I  �  =  M  '  %'  �   .�S  T?  �  f  {  '  $%  �  �   .�S  05  �  �  �  '  $%  �   .�S  $S:  �  �  �  '  �"  �   .�>  2hL  �  �  �  '  %'  �   .�>  CUB  �    $  '  $%  �  �   .�>  Q�2  �  =  M  '  $%  �   .�>  b�K  �  f  v  '  �"  �   .�4  qT  �  �  �  '  %'  �   .�4  ��K  �  �  �  '  $%  �  �   .�4  ��5  �  �  �  '  $%  �   .�4  �N.  �      '  �"  �   .U+  �)  P  8  H  '  �  �   .��  �!1  m   a  l  '  %'   .��  ��T  m   �  �  '  �  �  %'   .��  ��O  m   �  �  '  �  �  %'  �  �   .��  	;.  m   �  �  '  $%   .��  (	�B  m     $  '  �  �  $%   .��  C	�,  m   =  W  '  �  �  $%  �   a  1!T  �"  2�E    2�F  �   �&  �7  P  Qf Q� )�  3�~ 1�  4 }  4�} 4�} 4�� 4j| 4�| 4[| 4�} 4y| 4Dy 	4{ 
4_ 4Sy  5} C�   �  5�} F�  5�} L�  5�� O�  5m| R�  5�| U�  5^| X�  5�} [�  5|| a�  5Gy g�  	5{ l�  
5b r�  5Vy x�   6!| �0   &   &    )� ��  7!| �  �  H'  N'   8!|  �  �  H'  �   9ǁ $�         H'  m    ,� �� �     T'    �8 �  �� :	[ OB    �   ;<;   <�  =�  >�  ?;   =;   @int A�  <�  $   �/"  �  $,�  -�  K  :�!  �e  =�  � ?�$  "  @$%  �4  An%  �J  Bt%  �A  O�   �   z%   �A  Q!  !  z%  �%   �A  V*!  5!  z%  m    �
 Y51  �   M!  X!  �%  �    �
 ]�R  �   p!  {!  �%  �    � c?  �   �!  �!  z%  �   %   _ m.   �!  �!  z%  �   �    �3  q89  �   �!  �!  �%   B_Tp �"   �   ZD  8E  CU  A�&  "  Z'  m    D9+  N�&  Z'  m     A�  Ao  A�  A�  A�  A�  A�	  A(  A#  A�� A�� A�� 2*  7�"  E8   A�  �  /"  �  R"  �O 6"  �O Y"  pW   ="  qW  !m     "K"    #g"  ` &R"  ` '/"  �^ (Y"  �^ )6"  �T *m   �T +="  iY ,g"  hY -K"  �e 0R"  �e 1/"  [ 2m   [ 3="  Q 4m   Q 5="  �_ 6g"  �_ 7K"  �] :m   �] ;="  �Q >g"  �Q ?K"  .  <�"  `  Dm   �  W�"  �  _�"  �  em   t   mm   a  um     ~m   �  �m   3  �m   �  �m   H  �m   y  �m     �m   s  �m   T   �m   �  �m   F  �m   �  �m   �  �m     �m   V  �m   <�"  A�  s  N�"  �  V�"  \	  2m   o  7m   �  <m   �  Cm   �  m   <#%  F<*%  �"  GpO qO !/%  =   =P  <P  <   =w  AYe A�[ =�"  =*%  <�   =�!  <�!  <�  =6  A  �  8�&  �{  �$   ]�  �$  \�   �$  �D  !�$  �3  "�$  U>  #�$  &�  $�$  �  %�$  �*  &�$   ڡ  '�"  $�U  (�"  %TL  )�"  &�I  *�"  'Q  +�"  (�C  ,�"  )�J  -�"  *1  .�$  ,o(  /�"  0�U  0�"  1PL  1�"  2�I  2�"  3Q  3�"  4�C  4�"  5�J  5�"  6 H)%  K�$  �&  m   $%   IGT  P�&  <�%  �   m   m   <\  <�  <P  <a  =a  =�  ?P  =P  JD"  B'  K <W  <�  =+   <+   <�&  L�!  �'  MXF  AZ'  M\;  Am   NO�T  C�&    P  �'  �'  Qh  �'   '  L�  �'  NR__p �H     L"  �'  MXF  NZ'  M\;  Nm    P�  �'  (  Qh  (  S__a �(   '  �%  P�  (  2(  Qh  2(  Q#  '   H'  P�   E(  O(  Qh  O(   z%  P�  b(  l(  Qh  l(   �%  P!  (  �(  Qh  O(  Q#  '   P  �(  �(  Qh  l(  Q#  '   P�   �(  �(  Qh  O(  �(   �%  P  �(  �(  Qh  l(  S__a 	s�(   �%  P
  )  )  Qh  �'   PV  #)  -)  Qh  �'   T�  >)  Q)  Qh  Q)  Q#  '   '  P  d)  w)  Qh  w)  Q#  '   '  U(  ـ  �   ��)  �)  V(  � W/�X� �   U(   0�!   ��)  �)  V(  � Y(  8�   $�)  Z(  �( [D� \Q��1   P�   *   *  Qh  2(  M~  �   U�)  ԁ `��   �;*  ?,  V*  � V*  �]V)  ��p !?+  Zd)  �( ^)  ��� #�*  Z#)  �( _�'  ��   -Z�'  �(   `�'  ��� #Z�'  ) Z�'  1) a��   Z�'  O) Z�'  |) ]�'  ��� �3+  Z�'  �) Z�'  �) b`'  ��� VZu'  �) Zj'  �) c� d�'  �)    eʳ�     YV)  ϳ7   !+,  Vd)  ut�f)  ϳ   #�+  V#)  ut�_�'  ϳ   -V�'  ut�  _�'  ׳/   #V�'  us�Z�'  �) a�   Z�'  �) Z�'  $* ]�'  �� �,  g�'  Z�'  7* b`'  �� Vgu'  Zj'  7* c� h�'  S   e��     [}�[��e��1   iU  =K,   �#  i�   >K,  iB  ?K,  i�  Et,   �#  iB   Ft,  iC  Gt,  ie  Ht,  i8  It,  i�  Jt,  i

  X�,   �#  i�  Y�,  i�
  Z�,  j�   `�,  �#  i�  f�,   �#  i�  g�,  i�  h�,  i�  n$-   $  i�	  o$-  i�  p$-  iH  vM-   $  i`  wM-  iw  xM-  i   yM-  i~  �-   $  i   ��-  i�  ��-  i  ��-  i�   ��-  i�  ��-  i�	  ��-  i�  ��-   )$  i  ��-  i  ��-  i�  ��-  i�  �.   4$  i�  �.  i�  �.  i�  �.  im  �E.   ?$  i	  �E.  i2	  �E.  i�  �E.  i9  �E.  i[  ��.   J$  iJ  ��.  i�  ��.  i7  ��.  i�  ��.   U$  iI	  ��.  i$	  ��.  i�   ��.   `$  iN  ��.  ip  �/   k$  i�  �/  i:  �/  i�  �/  id   �/  i�  �B/   v$  i  �B/  i�  �B/  i�	  �k/   �$  i�  �k/  i  ؈/   �$  i�  و/  i�  ڈ/  i�  ۈ/  i+  �/   �$  i�  �/  i�   �/  i  ��/   �$  i�
  ��/  i�  ��/  i  �0   �$  i   �0  iF  �0  i�  �80   �$  i�  �80  i�  �80  iD  Oa0   �$  i�  Pa0  i1  Qa0  i�  W�0   �$  i^  X�0  i�  3�0   �$  i�  4�0  i�   8�0   �$  i�  9�0  il	  =�0  �$  iN  >�0  i^  ?�0  iL  @�0  ia  D1  %  iB  E1  i�	  F1  i  G1  i  H1  iy  I1  i�   c1   %  i�  !c1  k5   l�   l  l  l  l'  l3  l?  lK  lW  lc  	lo  
l{  l�  �  �1  �1  H    m>  Y  H     W   ��  �� 5� s� �     �i std  W	  %  0@�  �=  �  �b  ��	  Fe  �	  �3  �=  z   �  �   	J   
eq �<-  �  �   �  �   
lt ��1  �  �   �  �   ��  eF  �	  �   �  �     �K  �9    �   �   �(  
!  �    �    �   1  �A  �  ?  �  �     �5  �'  �  c  �  �     �3  �A  �  �  �    J    +  :  J   �  �   	U   �C   �P  U   �  �   �B  $6  �  �  �  �   eof (�:  U   ?  ,N0  U   �    _� ��	  �?  ��	  5�  6�  7  W  3�  �4  �$  q-  c=  o'  �5   �%  � �8  �X)  ��%  ��  �aO  �Y=  � P  �� �C  ��wS  ��O  � �?  ��5  �� 
$ g�  )W  �   �U  �A  �8  �P   EH  �� �4  �&  O   �7  (  �Q  G  �� ��  �M  �R   �-  �1  lO  �� b4 I  �9  i�  �N  �&  �  J�  �P  �1  �4  �  	}  dec �  t-  �  hex �  r'  �  < �   oct �  @� �  �[)  �   �%  "�   �  &�   dO  )�   \=  ,�   �P  /�    �C  3�   @zS  6�  ��O  9�  J�?  <�  �7  N�  	p  (  Q�  �Q  V�  O  Y�   app l�  	V  ate o�  in w�  out z�  �P  }�   beg �'   	c  cur �'  end �'   �Y  ,  �_ 
��  �M  
��   �_ 	.}  �  .  4  �   �  
��e  �  �  :    	R  Ic  ;�d  4  �  �  �  �   Fe  
?U   	�  {'  
E,  !T  �	  �E  >   Ic  
�A� E      �   &� 
GI   �M  ;  �* �e  �  N  T  �   �b  ��	  �* �_e  �  y    �   \b  (a  �  �  �  �   cb  �Pc  �  �  �  �	   �a  R(b  �  �  �  �   Fe  �U   �c  <�c  �    	  �   !a  *�a  �  "  (  �   !T  �	  �E  >    b�  c@  eK  fc  gx  h�  i�  j�  k�  l�  m  q*  rO  tn  u�  v�  x�  y�  |�  ~  �  �(  �B  �T  �j  ��  ��  ��  �>  b  �E  �  3F  ;�S  �  ,  2  �   9U  ؍0  p  J  P  �   �M  ��B  p  h  n  �    eU  ��4  �  �    p    bU  �IQ  �  �    p   !T  �	  �E  >   !�1  )�%  �    p    	
  	,  "�*  ��  �  �  �   "	W  �l  	  r  �   	�  "*  ��  7	  �  �   #�b  ��  $_Tp �	  �  �    %$   Ex	  �  $,  -   &�  &o  &�  &�  &�  &�  &�	  'int &(  &#  &�� &�� &�� %2*  7�	  (80    _� ԍ	  &�  �  x	  pW   �	  qW  !�	    "�	    #�	  )Fd 
  .  <
  `  D�	  �  W
  �  _
  �  e�	  t   m�	  a  u�	    ~�	  �  ��	  3  ��	  �  ��	  H  ��	  y  ��	    ��	  s  ��	  T   ȩ	  �  Щ	  F  ש	  �  �	  �  �	    �	  V  �	  *�	  &�  +s  N�	  �  V�	  \	  2�	  o  7�	  �  <�	  �  C�	  �  �	  *�	  	\  $
  gX  $
  X\  &�  X\  X,�  ,$Z  ./
   ,\ /�	  ,� 1�  ,Z  2�	  ,K]  3�	  ,�_  4�	  ,\W  5�	  ,�Z  6�	  ,-_  8�   ,VY  9  $,`  :'  (,�Y  ;<  ,,7_  <Q  0,BY  ={  4,b\  >Q  8,\  ?Q  <,7Y  @Q  @, Z  A�  D,SX  B�  H,n4 D
  L,`  F�  P,*5 G�  T -�  �  8  �	  �   *�  *�  -�      �	  �   *  .*�  -�	  '  �  �  �	   *  -�  <  �   *-  -�	  Q  �   *B  -�  p  p  p  �   *v  	�	  *W  /�  �   *�  0pO qO !�  1J   1z   &�  *z   *J   1�  &  �  8�  ,�{  +   ,]�  +  ,\�   +  ,�D  !+  ,�3  "+  ,U>  #+  ,&�  $+  ,�  %+  ,�*  &+   ,ڡ  '�	  $,�U  (�	  %,TL  )�	  &,�I  *�	  ',Q  +�	  (,�C  ,�	  ),�J  -�	  *,1  .+  ,,o(  /�	  0,�U  0�	  1,PL  1�	  2,�I  2�	  3,Q  3�	  4,�C  4�	  5,�J  5�	  6 ")%  K+    �	  p   2GT  P#  *�  	�	  *R  1I  *�  �^  !�  3Z  1]  ]   *�  "aY  ��	  x  ]   4\  C�	  �  ]   4xZ  M�	  �  ]   "`  ��	  �  ]   4�^  r�	  �  ]   4_X  ��	  �  ]  �   *@  4�_  �+    +  �	  ]   "�\  �]  *  p  p   44Z  ��	  O    �	  �	  ]   "7`  �]  n  p  p  ]   4>]  	�	  �  ]  �	  �	   4�Z  �	  �  ]  �   *�  	@  4�Y   �	  �  ]   4�Y  ��	  �  ]   5\  ��	  "�_  0+    +   3�]  W  p   "D[  T�	  (  p   "�[  a�	  B  p  p   3�\  )T  ]   6Y@ �j  ]  +   "�[  ©	  �  ]  +  �	  �	   2�]  i]  "D]  w+  �  +   4}W  ��	  �  �	  ]   *,  *�  7  �  �  8h  �   	�  *T  *�  75      8h     	�  7`  )  3  8h     7  A  W  8h  W  9__n �   	�  72  j  t  8h  �   7P  �  �  8h  �   7�  �  �  8h  W  9__n ��	   :�  �  9__c  �   	�  7�  �  �  8h  W  ;<�&  T�    7�       8h  W  ;<�&  >�    :�  ;  =hR  $;  =mR  $@   	�  	�  >�  :�  l  ?__a ��  ?__b ��   1	  1�  :�  �  ?__a ��  ?__b ��   	r  :	  �  ?__a ��  ?__b ��   7�  �  �  8h  �   	:  1)  :7	    $_Tp �	  ?__a �  ?__b �   	�  	�  *
  7n  *  ?  8h  ?  @�%  �p   	  7�  R  g  8h  ?  @�%  �p   7	  u  �  8h  W  ;<�&  ,�    *I  A�  �S  ��  �  Bh  �  � C__n <�  �D �  E�$  BR  �_D8 �  F�*  Ep  L* Dh   F�^  H�  �* F(  I�  �* G__c J�  �* FAc  M�  '+ H�  e�� J�  I�  �* Je�   �  K�  L�  n�   VI�  S+   M�   I�  f+ M�   K�     N� O�a  S�  Hg  t�� _�  Iu  y+ N� P  �+ Q�  v�  .P  I   y+ D  -  P
  �+ L�  }�   BR�  I�  �+   M͵   I   , M͵   K
     L�  ��4   /I�  !, J��   �  K�  L�  ��   VI�  4,   M��   I�  G, M��   K�       H3  ��8 X�  IA  Z, RJ   S�  ��P ZI�  m, NP K�  L�  ȴ   VI�  �,      HD  �h y�  I[  �, IR  �, Tx  �   ��  I�  �, I�  �, UK  �   �I`  �, IU  �,   VS�(   H  K�� {�  I3  - I*  '- TK  S�   ��  I`  - IU  :-  V`��   J�F   �  W�  HD  �� ur  I[  N- IR  n- Tx  �   �h  I�  N- I�  �- UK  �   �I`  N- IU  �-   V.�(   V�-  V@�@  VN�(   V��-  V �@  VZ�@   X>�Vµ    VI�K  Vc�K   	�  *�  %   �  Y�  	�  1�  ZU  =�   	9
  Z�   >�  ZB  ?�  Z�  E(   	D
  ZB   F(  ZC  G(  Ze  H(  Z8  I(  Z�  J(  Z

  Xu   	O
  Z�  Yu  Z�
  Zu  [�   `�  	Z
  Z�  f�   	e
  Z�  g�  Z�  h�  Z�  n�   	p
  Z�	  o�  Z�  p�  ZH  v   	{
  Z`  w  Zw  x  Z   y  Z~  6   	�
  Z   �6  Z�  �6  Z  �6  Z�   �6  Z�  �6  Z�	  �6  Z�  ��   	�
  Z  ��  Z  ��  Z�  ��  Z�  ��   	�
  Z�  ��  Z�  ��  Z�  ��  Zm  ��   	�
  Z	  ��  Z2	  ��  Z�  ��  Z9  ��  Z[  �:   	�
  ZJ  �:  Z�  �:  Z7  �:  Z�  �o   	�
  ZI	  �o  Z$	  �o  Z�   ��   	�
  ZN  ��  Zp  ��   	�
  Z�  ��  Z:  ��  Z�  µ  Zd   õ  Z�  ��   	�
  Z  ��  Z�  ��  Z�	  �   	�
  Z�  �  Z  �<   	�
  Z�  �<  Z�  �<  Z�  �<  Z+  �q   	�
  Z�  �q  Z�   �q  Z  �   	
  Z�
  �  Z�  �  Z  ��   	  Z   ��  ZF  ��  Z�  ��   	   Z�  ��  Z�  ��  ZD  O   	:  Z�  P  Z1  Q  Z�  W>   	E  Z^  X>  Z�  3[   	P  Z�  4[  Z�   8x   	[  Z�  9x  Zl	  =�  	f  ZN  >�  Z^  ?�  ZL  @�  Za  D�  	q  ZB  E�  Z�	  F�  Z  G�  Z  H�  Zy  I�  Z�      	|  Z�  !  \�  ]�  8  @  8   \�  1  ^>  Y  8    �   ��  c� � k  �     �n std  �   ��  ��   �   �    ��  �W   ]   �    W� 0   r   }   �   �    (� @� �   0   �   �     	�� 
0    0   int �   
�   �  �   ]   �   �   h  �   #  �    
�   
�   }   p�   �    h    �  
�   �   P� ��   �?  V  �   � ��� �   �   -� ��!   �q  �  �   � �   ��   �  �   �- �� ���   �  1  �  �       (�  � Q� k  �     �o �?  �0   (  �     �  r� g�   �� q}   �� � �� ��  �� j�   �� n0   	�� {ԇ �  �   �   
�   	� ą �  �   �   
�   �� �ˆ %   �   
�     �  	� �;  �  �� �� u� l� �� V� �  6� ��  � �(   �� ��   .� �/  �� ��  6� ��  
6  /    Ç �-  � �(   M� ��   $� ��   �� ��   Ŋ �/  Ç ��  �  
<  /   Ç �    
<  B   �  �Ȅ H  !  
<  B    �  �� �� �   J  d  
�  %   (  �  (   �� � � �  �   �  
�  �  (  �    �   I   �� �  �  �� !�  ˋ � W�  �    ��  N  �� N  �� U  ��   %  
l  r  /   �� �  :  E  
l  
/   �� O%� �  �  e  �  
�  %   �   �  (  �  (  H   �  Ɖ �   �  �  �  
�  %   (  �  (   �� 0� �  �  �  
�  �  (  �    �  ,�  ->   �� I�  /  T 0   (  %    �� I(  L   T (  %    F� R(  k  (  �  %    t� _�  �  �    �� g�  �  �    (� c�  �  �    !�� |�   *�  �   "�  �  "�  #abi �>   $std  (  �   U  x�� �    
      �  _� �7    ".  %&int ";  "�  '-  '�  �  (I   e  )e    �  "�  "x  }  �  "�  ';  "�  0   *  �  T 0   +WC  I(  +,� I%    */  �   T +WC  I(  +,� I%    ,%  �    -h    -#     l  /  "  '  ,�  ,  A  -h  A  +:� xF       ,�   Y  c  -h  c   �  ,�   v  �  -h  c   ,�   �  �  -h  c   *L  �  +� R(  +�� R�  +,� R%   ./`� V(    *k  �  +� _�    ,�  �  d  -h  d  +j� !%   +�� "(  +�� #�  +� $(  .0i )  ./WC  .(  /,� /%   /�� 0�  /,� 9�      �  ,2  w  �  -h  �  +j� �%   +�� �(  +�� ��  +� �(   �  ,�  �  �  -h  �  +�� �/   <  *�  �  +� g�    *�    +� c�    ,E    	  -h  d  +j� P%   +� Q�   +�� R�  +�� S(  +�� T�  +� U(  +�T  V	  1n� x./�� q(  /ۊ t�  /��  u�  /@� w�  .0i y  ./�� {�  /WC  |(  /T� }�   /,� ~%   /�� �  /g� ��  2�  /ӊ ��   ./�� ��   /�� ��        H  ,x  +	  >	  -h  >	  3d �/   6  ,�  Q	  �	  -h  d  4dst 1�  5�� 1(  5�T  2�	  .6.� 7/  .7i ;  .6�� =;  6WC  >(  6,� ?%   6�� @�  6�� A�      �  8�  a� ��   ��	  
  9�  � :϶;� �   8�  �� ж!   �)
  ]
  9�  � <�  ض   S
  =�  �- >� ?��   @�  Ɖ  ��   �x
  �  9�  � 9�  �9	  �9  �9  �A  ��� &�
  =,   . =5  . B��   C  =  H. =  h. =	  �. =�  �. =�  �. C D+  �. C0 D5  2/ E@  PFK  DV  `/ <�  7�   /O  =�  ~/  G�  H�H 7=�  �/ =�  �/ =�  �/ HL�   �  D�  
0 I�  L�   X=�  0 =�  
0   I�  W�   [=�  A0 =�  T0       @  %� �o  ��  �  9  � 9  �9(  �93  �9>  �9I  �9T  �9_  �Jj  K` �  Fr  F}  F�  F�  I  7�-   [=,  r0 =5  �0 BR�    C� =_  �0 =T  -1 =I  Y1 =>  �1 =3  �1 =(  �1 =  	2 =  52 C� Lj  }�C� Dr  l2 D}  �2 D�  !3 D�  �3 A  '�� b5  =,  =4 =5  i4 B>�   K� �  D�  �4 C E�  �LD�  �4 D�   5 E�  PF�  D�  J5 KH �  D�  �5 D	  �6 Ai  ��x �4  =�  �7 =�  �7 =�  28 =�  �8 =w  �8 A�  ��� ��  =�  )9 =�  w9  M��A   =�  �9 =�  �9 =�  �9 =�  �9 =w  	:   Gi  �� �=�  : =�  I: =�  u: =�  �: =w  ; <�  ��   ��  =�  0; =�  [;  M��6   =�  �; =�  �; =�  �; =�  �; =w  �;    A�  �� {�  =�  �; =�  <  <�  �   ~  =�  w<  A�  �� ��  =�  �< =�  �< =�  = K u  D�  %= G�  �0 X=�  := =�  %=   I�  .�   [=�  \= =�  o=   CH D�  �=    I�  ��   g=�  �= =�  �=      @C	  � `�Q  ��  �  9Q	  � 9Z	  �9f	  �9r	  �Hg�"   &  F	  B|�d   C` =r	  > =f	  2> =Z	  R> =Q	  r> C` D	  �> C� D�	  �> C� E�	  �PD�	  T? E�	  PF�	  F�	  N�  ��   ?�  =�  ?  N�  þ   H;  =�  �? =�  �? =�  �? HǾ     D�  �? I�  Ǿ   X=�  @ =�  �?   I�  Ͼ   [=�  *@ =�  =@   N�  �   NY  =�  Q@  N	  X�#   =�  =4	  e@ =+	  �@  Oh  {�� A�  =v  A  OK  }�� @�  =Y  ?  P  �+   w=,  SA =5  gA B/�        Q�  R�  1       STmw  ww  /  r  r    v    ��  � �� k  (     �s std  �e  Ӫ  ��   �f   ptr f   � ��h   � �   �  �1  	f     �   �  � Ԍ k  8     {t �  (  _� �>   �  �  P   �  �  o  �	  �  qW  !~   int   "�   �  #  s  NE   �  VE   .  <s   `  D~   �  Ws   �  _�   �  e~   t   m~   a  u~     ~~   �  �~   3  �~   �  �~   H  �~   y  �~     �~   s  �~   T   �~   �  �~   F  �~   �  �~   �  �~     �~   V  �~   %   �  \	  2~   o  7~   �  <~   �  C~   �  ~   *    �  ~    	rem ~    +   �  #@  A  �  $,    	rem %,    A  &  
std  �  	v  	wA  	{�  	�  	�B  	�W  	�l  	��  	��  	��  	�  	�  	�I  	�i  	��  	��  	��  	��  	��  	�  � �� 
Z  �� 
W   � �~          �  >0  0  7   �� =  %   �  H~   W  7   �  I,   l  7   �  �   �  �  �  3   3   �   �  �  ~   �  �  �   div   �  ~   ~        ��  �  7   �   A    ,   ,    �  .~     7  3    �  \3   <  <  7  3    B    3  >~   i  <  7  3    �  �  �   3   3   �   k� q~   �  |�  l      W0  �  7  �   �    f,   �  7  �  ~    �  g>     7  �  ~    ?  �~     7      %  A  P>�  �  A   t  B  +  F�  �  G�  �  J"  p  N~   p  Y~     Z(  �  [(   �  \C  $w  ]�   (4  a�  0 �  ��  �  �"   �  �l    �  �:  �  �:  P  @�   ++CCUNG}  L�  ++CCUNG �  abi �  + 0l   (  5l   �  =�   B�  �  �   �  M  3  �  ]  K  	  �   �  LY  �  W�  �  �  �  �   �  ^   Z  �  \N   �  ]�  V  b8  `  c8   �    �      $  .  P   *  �   �  ��   � �  ��   �!D  Oj   �   !�  Pj  !1  Qj  !�  W�   �   !^  X�  !U  =�   �   !�   >�  !B  ?�  !�  E�   �   !B   F�  !C  G�  !e  H�  !8  I�  !�  J�  !

  X&   �   !�  Y&  !�
  Z&  "�   `O  �   !�  f`   �   !�  g`  !�  h`  !�  n�   �   !�	  o�  !�  p�  !H  v�   �   !`  w�  !w  x�  !   y�  !~  �     !   ��  !�  ��  !  ��  !�   ��  !�  ��  !�	  ��  !�  �@	     !  �@	  !  �@	  !�  �@	  !�  �u	     !�  �u	  !�  �u	  !�  �u	  !m  ��	   $  !	  ��	  !2	  ��	  !�  ��	  !9  ��	  ![  ��	   /  !J  ��	  !�  ��	  !7  ��	  !�  � 
   :  !I	  � 
  !$	  � 
  !�   �I
   E  !N  �I
  !p  �f
   P  !�  �f
  !:  �f
  !�  �f
  !d   �f
  !�  ɧ
   [  !  ʧ
  !�  ˧
  !�	  ��
   f  !�  ��
  !  ��
   q  !�  ��
  !�  ��
  !�  ��
  !+  �"   |  !�  �"  !�   �"  !  �K   �  !�
  �K  !�  �K  !  �t   �  !   �t  !F  �t  !�  �   �  !�  ��  !�  ��  !�  3�   �  !�  4�  !�   8�   �  !�  9�  !l	  =   �  !N  >   !^  ?   !L  @   !a  D5  �  !B  E5  !�	  F5  !  G5  !  H5  !y  I5  !�   �   �  !�  !�  #�  D�  FN  $�   ++CCUNG$  ++CCUNG \   ��  �� �� k  �     �v �  (  _� �>   �  �  P   �  �  o  �	  �  qW  !~   int   "�   �  #  s  NE   �  VE   .  <s   `  D~   �  Ws   �  _�   �  e~   t   m~   a  u~     ~~   �  �~   3  �~   �  �~   H  �~   y  �~     �~   s  �~   T   �~   �  �~   F  �~   �  �~   �  �~     �~   V  �~   %   �  \	  2~   o  7~   �  <~   �  C~   �  ~   	*    �  	~    	rem 	~    +  	 �  	#@  A  �  	$,    	rem 	%,    A  	&  
std    
v  
wA  
{  
�5  
�\  
�q  
��  
��  
��  
�   
�  
�6  
�c  
��  
��  
��  
��  
��  
��  
�  � �� Z.  �� W.  z0  �]A  �  �  f.   � 	�~   .  .   4  �  	>J  J  Q   �� W  %   �  	H~   q  Q   �  	I,   �  Q   �  	�   �  �  �  3   3   �   �  �  ~   �  �  �   div 	  �  ~   ~        	��     Q   �  	 A    ,   ,    �  	.~   6  Q  3    �  	\3   V  V  Q  3    \    3  	>~   �  V  Q  3    �  	�  �   3   3   �   k� 	q~   �  	|�  l      	WJ  �  Q  �   �    	f,   �  Q  �  ~    �  	g>     Q  �  ~    ?  	�~   3  Q   + 0l   (  5l   �  =�   B�  �  �   �  M  3  �  ]  K  	  �   �  LT  �  W�  �  �  �  �   �  ^   Z  �  \I   �  ]�  V  b3  `  c3      �  A  P>�  �  A�   t  B�  +  F�  �  G�  �  J�  p  N~   p  Y~     Z�  �  [�   �  \>  $w  ]�   (4  a�  0 �  ��  �  ��   �  �l    �  ԰  �  �    �� t�   �  �    �  W�    I   �� �   )  �    �  (�   >  �    !�  ^"P  @3   ++CCUNG"}  L3  ++CCUNG#�  XC	  #�  [C	   �  $abi �  �  �  �    �    �  P   %  &�  �  'exc ��   &�    (eo t�  )*e  w�    &�    (c WI   +  ��   �Q  ,0  �   � -��   .�� !�  �   +)   �~   �C	  ,0  (�   � /P 0�� *�  ~A 0�  ,C	  �A 0`  -�  �A 1e  .�  1�� /�   0�� B~   �A 2  �p 5�  3  ?B  4�  �   .	  3�  lB  4�  Z�   R/	  3�  �B -Z�   5�    6�m  6~�    �  +>  ��|   ��	  /� 0�  `C	  �B 0e  a�  �B 0�� q~   
C 4  ��   j�	  3  hC  6��y  6��R  6��    +�   �   ��	  -�   0�  �C	  �C 6�m    7D  O

   �   7�  P

  71  Q

  7�  W3
   �   7^  X3
  7U  =P
   �   7�   >P
  7B  ?P
  7�  Ey
   �   7B   Fy
  7C  Gy
  7e  Hy
  78  Iy
  7�  Jy
  7

  X�
   �   7�  Y�
  7�
  Z�
  8�   `�
  �   7�  f    �   7�  g   7�  h   7�  n)   �   7�	  o)  7�  p)  7H  vR   �   7`  wR  7w  xR  7   yR  7~  �     7   ��  7�  ��  7  ��  7�   ��  7�  ��  7�	  ��  7�  ��     7  ��  7  ��  7�  ��  7�  �     7�  �  7�  �  7�  �  7m  �J   $  7	  �J  72	  �J  7�  �J  79  �J  7[  ��   /  7J  ��  7�  ��  77  ��  7�  ��   :  7I	  ��  7$	  ��  7�   ��   E  7N  ��  7p  �   P  7�  �  7:  �  7�  �  7d   �  7�  �G   [  7  �G  7�  �G  7�	  �p   f  7�  �p  7  ؍   q  7�  ٍ  7�  ڍ  7�  ۍ  7+  ��   |  7�  ��  7�   ��  7  ��   �  7�
  ��  7�  ��  7  �   �  7   �  7F  �  7�  �=   �  7�  �=  7�  �=  7�  3f   �  7�  4f  7�   8�   �  7�  9�  7l	  =�  �  7N  >�  7^  ?�  7L  @�  7a  D�  �  7B  E�  7�	  F�  7  G�  7  H�  7y  I�  7�   "   �  7�  !"  I  9E   ++CCUNG9Y  ++CCUNG:�� ��    �   ��  i� ,� k  �     ;y (  �     �   "� �>   �   �    6� #>   n   y   "     K� ��� >   �   "    	� 0�   �    "� !�   �   �   (     
K� 5֎ �   �   (     �  abi �3        int   �5     >   �   std  A  �z I�  �  �   �z L`  f  A   � 9  {  �  A     (� /c� G  9  �  Y    �� <�  6  ��    �� �  �  _  e   �� ?�  �  _   X� �      _     (� &�� G  �  /  k    9  �   9  M  R  �  6  �  ;  ;  �    �  h  �  #  �   _    f  �  �  h  �  #  �   A    �   �  �  h  �  #  �   (    Z        h    #     "    q  X�  �   �8  A    �  �  l� 0�   �\  e  �  �    @�   �|  �   h  �  �  k  �  P�   ��  �   h  �  �  Y  q  � `�   ��  �    � !e��  "� �   �  �� p�   �  #  �  � !u��  "� �   �  � ��   �>  G  �  �  �  3� ��   �b  }  �  � !���  "� �   �  �� ��   ��  �     �  �  �� ��   ��  �     � !���  "� �   #�  1  �  �   $ �   ��  � �� k  @     �z (  �     �    >   �� o   �� !ˋ � W�   	�   
,�   
-3   �� |�   
*o    C   �  abi �3   std  �  � X�   �  � �   F�  ��  �� �   �     �  �   H�  cÑ �    !  �   �3 s�� �   9  D  �  �   U  x�� �   \  g  �  �   2  �ܓ �     �  �  �   �� 7�� �   �   �  �  �   p� >� �   �   �  �  �   :� E�� �   �   �    �  �  �  �   �� LE� �   �   +  ;  �  �   �   � �K  V  �  �   �  �ۑ �  m  x  �  �   � ��  �  �    �    int �  �   �  �5  �  �  �  �  �   �  �  �  �  �    �   �    !h    !#     �  �   D  )  >  !h  >  ":� xC   �  �  #�  &� ��   �c  l  $�  �  %�  ��   ��  �  &h  >  �  %�  ��   ��  �  &h  >  �  %  ��   ��  �  &h  >  � '�   �'�  � #�  Ӓ  �   �    $�  � (��  )� �   %�  �I   �5  �  &h  >  � *�� F�  �'�  �'�  �+  !�( H$)  � ,2  �C -6��    �   .�   /�  1  �  �   0mw  ww  �  �  �    
   w�  �� Ԕ k        )| �?  �0   (  �     q  r� g�   �� q}   �� � �� ��  �� jq   �� n0   	�� {ԇ w  �   �   
~   	� ą w  �   �   
~   �� �ˆ %   �   
~     ��    	� �C  �  �� �� u� l� �� V� �  6� ��  � ��   �� �  .� ��  �� �q  6� ��  
�  �    Ç �5  � ��   M� �  $� �  �� �  Ŋ ��  Ç ��  �  
�  �   Ç �
    
�  �   �  �Ȅ �  )  
�  �    �  �    O  Z  
�  �   �  1� �  p  {  
�  �    ��  �  
�     �� �   �  �  
�  
�   �� -�� w  �   �  �  
q  q     :�  � w  �       
q      "   �� ` � w  �   <  Q  
q  q  �  )   �� ��   i  �  
q  %   �  q  �   �� F�� w  �   �  �  
q  %     q  �  q  �  �   � :\�   �   �  
q  %   �  q  �    �   I   �� 4  �� !ˋ � W�   i   ,�   ->   !� kw  \     "�� |�    *4   #  �  #  $abi �>   %std  �  � �  U  x�� w  �  
  Z    �   #�  &'int #C  #�  (5  (�  #�   (  (�   #    �  #  )#�  �  (C  *�  =  P  +h  P  +#  U   �  �  (�  *�  n  �  +h  �  ,:� x�     Z  *�  �  �  +h  �  ,�� !  ,]� "  ,W� #"   q  *�  �  *  +h  �  %   ,� H  ,�� Iq  ,�� J�  ,�� Kq  ,� L�  ,�T  M*   �  *�  =  P  +h  P  -d ��   �  .G  k  ,� k   /�  `�X   ��  �  0h  �  � 1�� .q  �1�� /  �2l�G   3�T  1C  �`4/  l�   1�  5F  6=  �C  7U  ��x 48_  �d   9�  ��   �  N  0h  �  � :%   �1�� <�  �:q  �1� >�  � ;/  �� ��   �i  �  8=  � <��=� �   ;/  e� ��!   ��  �  8=  � 4/  ��   �  6=  -D >� ?��	   9   �a   ��  G  0h  �  � @dst aq  �@obj a�  �1�T  bG  �7`  7�� d8n  � 6w  LD AL��	    )  B�  � ��z   �g  �  8�  � 8�  �8�  �8�  �4`  ��   %�  6n  kD 6w  �D A���	   C� 6�  E 6�  $E 6�  CE 6�  bE   ;�  �� ��   ��  �	  8�  � 8�  �8�  �8�  �8�  �8  �8  �8  �D� �	  6�  �E 6  �E 6  �E 6  F 6�  1F 6�  fF 6�  �F 6�  �F 7`  -�� V6n  �F 6w  !G A@��	    E`  W�!   O6n  MG 6w  mG Aj��	    F\  G�  1  �	     Hmw  ww  �        �   ��  ֖ {� k  @     4~ std  �   z 6�   �   �    z U   `   �   �    z 9p   v   �    	�� 0   �   �   �   �    
(� c� �   0   �   �     �� 0    0   �   int �   �   �  �   v   �     h    #     �   �   �   ��   �1  >  h  >  �  �   �   �� ��   �^  u  �   � ��� �   �    ��!   ��  �  �   � �   ��   �  �   �G �� ��   �  �1  �  �    �   4�  � �� k  `     �~ std    v  6�  x  K�  �  M   x  Ob   m        	�  Qw  �   �      	�  R  �   �      
  T8    �   �   
   x  Z�   �      x  \�   �        x  _�       �   x  c  #       �  p�  !  ;  F       �  t�  !  ^  i       �  {y  �    '   n	 ~%  �  �    !   �  ��  .  �  �  
   �  �h  5  �  
    ;    :;   �  �  � �  vY  w�  {�  ��  ��  ��  �  �K  �f  �{  ��  ��  ��  ��  �  �*  �;  �[  �z  ��  3�  �� Z�  �� W�    X�  /  s�  �  7.  �  D  ֘ Jϗ �  �  �   � e� �  �    ;   �  �  �  ;   ;   int �  �  �  (  _� �T  �  �  �   �  ��    �  ��   #  �� !
  �[  �  �  �  �  o  �	  �  qW  !'    "�  �  s  	N�  �  	V�  .  
<�  `  
D'  �  
W�  �  
_�  �  
e'  t   
m'  a  
u'    
~'  �  
�'  3  
�'  �  
�'  H  
�'  y  
�'    
�'  s  
�'  T   
�'  �  
�'  F  
�'  �  
�'  �  
�'    
�'  V  
�'  ;  �  \	  2'  o  7'  �  <'  �  C'  �  '  "*  Y  �  '   #rem '   +   4  "#@  �  �  $B   #rem %B   A  &d  $� �'  �  �   �  %$�  >�  �  �   �� �  ;  $�  H'  �  �   $�  IB    �   $�  �  *  *  *  I  I  1   0  &7  ''  K  *  *   (div Y  f  '  '   $    ��  {  �   )�   �  �  B  B   )�  .'  �  �  I   )�  \I  �  �  �  I   �    )3  >'  �  �  �  I   *�      I  I  1   k� q'  +�  |;  �   $  W�  U  �  U   �  $  fB  z  �  U  '   $�  gT  �  �  U  '   $?  �'  �  �   �  =�     5  ,�  +:  �  �   ,�  =�  �  �   -�� �4� �  -�� �� �  .P  @~   ++CCUNG.}  L~  ++CCUNG /abi ��  0(�  1�  `  23ʗ Z�    1�  x  23ʗ u�    4�  �?   ��  5 +�  � 6��  6'��  6/��  68��  6F��  6O��   7�  P�   �	  8H  S�   9
	  9S�   :S  �G   6^�x   4�  `�   �?	  5 =�  � 6l��   7�  p�   ��	  8`  s�   Fy	  9s�   :k  �G   6~�	   7�  ��   ��	  ;ʗ J�  �G 9��
   <old L�  P  =H  �  ��   ��	  9��   >S  P  7�  ��   � 
  ;ʗ e�  �G 9��
   <old g�  P  =`    ��   �I
  9��   >k  P  ?D  	OU
   �  ?�  	PU
  ?1  	QU
  ?�  	W~
   �  ?^  	X~
  ?U  
=�
   �  ?�   
>�
  ?B  
?�
  ?�  
E�
   	  ?B   
F�
  ?C  
G�
  ?e  
H�
  ?8  
I�
  ?�  
J�
  ?

  
X     ?�  
Y  ?�
  
Z  @�   
`:    ?�  
fK   *  ?�  
gK  ?�  
hK  ?�  
nt   5  ?�	  
ot  ?�  
pt  ?H  
v�   @  ?`  
w�  ?w  
x�  ?   
y�  ?~  
�   K  ?   
��  ?�  
��  ?  
��  ?�   
��  ?�  
��  ?�	  
��  ?�  
�+   V  ?  
�+  ?  
�+  ?�  
�+  ?�  
�`   a  ?�  
�`  ?�  
�`  ?�  
�`  ?m  
��   l  ?	  
��  ?2	  
��  ?�  
��  ?9  
��  ?[  
��   w  ?J  
��  ?�  
��  ?7  
��  ?�  
�   �  ?I	  
�  ?$	  
�  ?�   
�4   �  ?N  
�4  ?p  
�Q   �  ?�  
�Q  ?:  
�Q  ?�  
�Q  ?d   
�Q  ?�  
ɒ   �  ?  
ʒ  ?�  
˒  ?�	  
ѻ   �  ?�  
һ  ?  
��   �  ?�  
��  ?�  
��  ?�  
��  ?+  
�   �  ?�  
�  ?�   
�  ?  
�6   �  ?�
  
�6  ?�  
�6  ?  
�_   �  ?   
�_  ?F  
�_  ?�  
�   �  ?�  
�  ?�  
��  ?�  3�   �  ?�  4�  ?�   8�     ?�  9�  ?l	  =�    ?N  >�  ?^  ?�  ?L  @�  ?a  D     ?B  E   ?�	  F   ?  G   ?  H   ?y  I   ?�   m   )  ?�  !m  �  A   ++CCUNGA   ++CCUNGBf� �C�    �     D�  E>  Y  �     F      �   *�  l� C� k  �     -� (  �  #  �� �  std  8  v  6  x  K�  �  M8   x  O�   �   	:  
8   �  Qw  �   �   	:   �  R  �   �   	:     T8  8  �   �   	@   x  Z�   �   	:   x  \    	:  
F   x  _  )  	:  

   x  c9  D  	:  
L   �  p�  R  \  g  	:  
F   �  t�  R    �  	:  
L   �  {�  �  	:  	X   n	 ~%  �  �  	:  
R   �  ��  _  �  �  	@   �  �h  f  �  	@    \    :\   �  �A   �   �� �� ?0  	�     \   �  �  \   \   int �       �  -� �X  �  
�   � .3   )� ȭ  
�  
X   q= �X  �  
�   
� � e= �X  �  
�   !Z� Q�  
�   "Y< x
�    #abi �l  $   �d  $*; 15  %�8  %�; %N;  &�� R  '�� �K  	�    (�= 5^      �  o  �  �  �  �	  �� �� �    )$  �  �  *h  �   �  5  )>  �  �  *h  �   �  �  +w    ,g ��   +�     ,g ��  ,v �X   +�  4  ,g ��   -�  .�  ��I   ��  /g ��  � 0   ��� M1*  H 2  ��   �  1  _H 1  sH  34  ��#   �2�  ��   ��  1�  �H  4��_  4	�r     .�  �	   �  5g Q�  � 6  �	   n7   8  �   .�   �   �Y  5g x�  � 6  $�   �7   8  �   9R   :�  8  r  
,    ;�  �  
8  
8  
�   �  <
8    /   p�  k� 2� k        h� �  �  (  _� �E   �  �  W   �  �  o  �	  qW  !~   int   "�   �  #  s  NL   �  VL   .  <s   `  D~   �  Ws   �  _�   �  e~   t   m~   a  u~     ~~   �  �~   3  �~   �  �~   H  �~   y  �~     �~   s  �~   T   �~   �  �~   F  �~   �  �~   �  �~     �~   V  �~   ,   �  \	  2~   o  7~   �  <~   �  C~   �  ~   *    �  ~    	rem ~    +   �  #@  A  �  $3    	rem %3    A  &  
std  1  	v  	wA  	{1  	�M  	�t  	��  	��  	��  	�  	�  	�3  	�N  	�{  	��  	��  	��  	��  	��  	�  	�6  
RK  
Ue  
[z  
\�  � �� ZF  �� WF  _� �E   �  f.   � �~   F  F   L  �  >b  b  i   �� o  ,   �  H~   �  i   �  I3   �  i   �  �   �  �  �  :   :   �   �  �  ~   �  �  �   div     ~   ~        ��    i   �   A  3  3   3    �  .~   N  i  :    �  \:   n  n  i  :    t    3  >~   �  n  i  :    �  �  �   :   :   �   k� q~   �  |�  %      Wb  �  i  �   �    f3     i  �  ~    �  gE   6  i  �  ~    ?  �~   K  i   ��  E~   e  i  i   ��  U�  z  ~    ��  O�  �  �  i   ��  F:   �  �  i  :    + 0%   (  5%   �  =�   B�    �   �  M  3  �  ]  K  	  �   �  L�  �  W-  3  C    C   I  ^   Z�  �  \�   �  ]"  V  b�  `  c�      6  A  P>.  �  AI   t  BZ  +  F  �  G  �  J`  p  N~   p  Y~     Zf  �  [f   �  \�  $w  ]�   (4  aI  0 =  Pp�    s�    �  xZ  +  |  �  }  �  �`  p  �~   p  �~     �f  �  �f   �  ��  $w  ��   (4  �I  0 �  d�   �       ��  �    Ϛ �H  � �  H   P  @�   ++CCUNG}  L�  ++CCUNG �  abi ��  �  Z  �    O  �  l  W   ��  !~   $   �
   *; 1�  �8  �; N;  !�; v_	  �= |q   "�; �  �  #
  "
   $�  ��= (
  �  �  #
  "
   %�; �
	  	  #
   &\ ��: $	  *	  #
   &f ��8 >	  D	  #
   '�9 ��: .
  X	  #
    �  !(8 ��	  (r< �  �9 �4
   "(8 �	  �	  #?
  E
   $�  �< K
  �	  �	  #?
  E
   )(8 ��	  �	  #?
  9
   *'8 ��	  #?
  #~     d	  +�= 5
   �   �� �� �  ,_	  ,�  q  9
  ,p	  d	  ,�	  ,d	  -2�  y� L%   .t
  /�� `�   -^c
  0�  �
  �
  1h  �
   
  2^�  �
  3w  �~   3-�  �~    0	  �
  �
  1h  �
   0*	  �
  �
  1h  �
   0�	  �
    1h    3F�  �   ?
  9
  0�	  $  7  1h    1#  7   ~   4�  0�z   ��  5Ú d  �H 6V  ~7� 8ret f�   �H 9`�J   �  :�_ md	  ;�� oX
  I ;��  p%   HI <��%   <B�    4�  ��<   �C  5�� ��   �I =��8   >WC  ��  �G�8ptr ��  �I 9��   8  ;��  �C  �I :�_ �d	   ?��%    %   .  4�  ��m   ��  6V  �7 8ret �H  %J 9 �=   �  :�_ �d	  ;�� �X
  eJ ;��  �%   �J <=�%   <��    4�  `�I   �F  5�� �H  �J =d�E   >WC  ƨ  @F�8ptr Ǩ  �J 9r�   ;  ;��  �C  K :�_ �d	   ?��%    @D  OR   �   @�  PR  @1  QR  @�  W{   �   @^  X{  @U  =�   �   @�   >�  @B  ?�  @�  E�   �   @B   F�  @C  G�  @e  H�  @8  I�  @�  J�  @

  X   �   @�  Y  @�
  Z  A�   `7  �   @�  fH   �   @�  gH  @�  hH  @�  nq   �   @�	  oq  @�  pq  @H  v�   �   @`  w�  @w  x�  @   y�  @~  �     @   ��  @�  ��  @  ��  @�   ��  @�  ��  @�	  ��  @�  �(     @  �(  @  �(  @�  �(  @�  �]     @�  �]  @�  �]  @�  �]  @m  ��   $  @	  ��  @2	  ��  @�  ��  @9  ��  @[  ��   /  @J  ��  @�  ��  @7  ��  @�  �   :  @I	  �  @$	  �  @�   �1   E  @N  �1  @p  �N   P  @�  �N  @:  �N  @�  �N  @d   �N  @�  ɏ   [  @  ʏ  @�  ˏ  @�	  Ѹ   f  @�  Ҹ  @  ��   q  @�  ��  @�  ��  @�  ��  @+  �
   |  @�  �
  @�   �
  @  �3   �  @�
  �3  @�  �3  @  �\   �  @   �\  @F  �\  @�  �   �  @�  �  @�  ��  @�  3�   �  @�  4�  @�   8�   �  @�  9�  @l	  =�  �  @N  >�  @^  ?�  @L  @�  @a  D  �  @B  E  @�	  F  @  G  @  H  @y  I  @�   j   �  @�  !j  B,   �  C�  D�  � >�� W{  �G>� XX
  �GB.  �  C�   > � Z�  @F>�� [X
  FEh
  F�	   �  G   ++CCUNGG!  ++CCUNG�� E�   %  :    H  ;�     �   1�  U� � k  �     · �  (  _� �>   �  #  �� �  �  c   �  �  o  �	  �  qW  !�   int   "�   �  s  NX   �  VX   .  <�   `  D�   �  W�   �  _�   �  e�   t   m�   a  u�     ~�   �  ��   3  ��   �  ��   H  ��   y  ��     ��   s  ��   T   ȑ   �  Б   F  ב   �  ��   �  �     �   V  �   %   �  \	  2�   o  7�   �  <�   �  C�   �  �   	*    	�  	�    
rem 	�    +  	 �  	#@  M  	�  	$,    
rem 	%,    A  	&(  std    
v  
wM  
{  
�7  
�^  
�s  
��  
��  
��  
�  
�  
�8  
�e  
��  
��  
��  
��  
��  
�  
�   v  6�  x  K�  	�  M�    x  O!  ,  5  �    �  Qw  ?  E  5   �  R  X  ^  5     T8  �   u  {  ;   x  Z�  �  5   x  \�  �  5  A   x  _�  �  5  �   x  c�  �  5  G   �  p�  M  �    5  A   �  t�  M    (  5  G   �  {8  C  5  �    n	 ~%  W  b  5  M   �  ��  S  z  �  ;   �  �h  Z  �  ;    �   :�  �  �S   � �  �� i0  z �  z 9�  �    ��    �� ?�  n    _� �>   �� q� �   � 	��   0  0   6  �  	>L  L  S   �� Y  %   �  	H�   s  S   �  	I,   �  S   �  	�   �  �  �  3   3   �   �   �  !�   �  �  �   "div 	  �  �   �        	��    S   #�  	 M    ,   ,    #�  	.�   8  S  3    #�  	\3   X  X  S  3    ^    #3  	>�   �  X  S  3    $�  	�  �   3   3   �   %k� 	q�   &�  	|�        	WL  �  S  �   �    	f,     S  �  �    �  	g>      S  �  �    ?  	ґ   5  S   �  �  '�  (�  '�  �  �  �   �  �  )�  �  �  *h  �   n  �  )�  �  �  *h  �   �  +�  *�  �   ��c   �M  ,sz *   3K -H .p ,�   vK /h B  0 4�  �K 1�  ��   6&  2�  �K  3��  3���  3��   3���    4D  OY   �   4�  PY  41  QY  4�  W�   �   4^  X�  4U  =�   �   4�   >�  4B  ?�  4�  E�   �   4B   F�  4C  G�  4e  H�  48  I�  4�  J�  4

  X	   �   4�  Y	  4�
  Z	  5�   `>	  �   4�  fO	   �   4�  gO	  4�  hO	  4�  nx	   �   4�	  ox	  4�  px	  4H  v�	     4`  w�	  4w  x�	  4   y�	  4~  �	     4   ��	  4�  ��	  4  ��	  4�   ��	  4�  ��	  4�	  ��	  4�  �/
     4  �/
  4  �/
  4�  �/
  4�  �d
   %  4�  �d
  4�  �d
  4�  �d
  4m  ��
   0  4	  ��
  42	  ��
  4�  ��
  49  ��
  4[  ��
   ;  4J  ��
  4�  ��
  47  ��
  4�  �   F  4I	  �  4$	  �  4�   �8   Q  4N  �8  4p  �U   \  4�  �U  4:  �U  4�  �U  4d   �U  4�  ɖ   g  4  ʖ  4�  ˖  4�	  ѿ   r  4�  ҿ  4  ��   }  4�  ��  4�  ��  4�  ��  4+  �   �  4�  �  4�   �  4  �:   �  4�
  �:  4�  �:  4  �c   �  4   �c  4F  �c  4�  �   �  4�  �  4�  ��  4�  3�   �  4�  4�  4�   8�   �  4�  9�  4l	  =�  �  4N  >�  4^  ?�  4L  @�  4a  D$  �  4B  E$  4�	  F$  4  G$  4  H$  4y  I$  4�   q   �  4�  !q  6�  �   �  >    7�  �  �   �   �   �  8�  �    9�� E�   3     �   f�  =� � k  �     �� std  �   v� ̠   �   �    v� �W   ]   �    � 0   r   }   �   �    (� � �   0   �   �     	�� 
0    0   int �   
�   �  �   ]   �   �   h  �   #  �    
�   
�   }    �   �    h    �  
�   �   � 0�   �?  V  �   � ?�� �   �   ˝ @�!   �q  �  �   � �   H�   �  �   �K T� a��   �  1  �  �    }   ��  C� � k  �     n� (  �     �  abi �3   $   ��   �� ��   �    �� �}   �   	�    
�� X   �   	�   	�      std  �   ��  X   int �   �   �   h  �   #  �    �   �   �   � p�   �    �   � �� �   �   Ҟ ��!   �7  k  �   � �   ��   a  �   �K �� ��k   �  1  ~  ~    0   I�  8� �� k  �     L� (  _� �7   �     �   �� /� 6P  @�   ++CCUNG}  L�  ++CCUNG �  abi �>   �  int �  =�   �  	std  �   
�  f.   �  �  �  �   �  o  �	  qW  !�     "�     #  #  s  N�   �  V�   .  <�   `  D�   �  W�   �  _  �  e�   t   m�   a  u�     ~�   �  ��   3  ��   �  ��   H  ��   y  ��     ��   s  ��   T   Ț   �  К   F  ך   �  ��   �  �     �   V  �   �  \	  2�   o  7�   �  <�   �  C�   �  	�   gX  
  w  I   ��   ��  ��  ���    P   ��   ��  ��  ���    D  O�      �  P�  1  Q�  �  W�   +  ^  X�  U  =   6  �   >  B  ?  �  E?   A  B   F?  C  G?  e  H?  8  I?  �  J?  

  X�   L  �  Y�  �
  Z�  �   `�  W  �  f�   b  �  g�  �  h�  �  n�   m  �	  o�  �  p�  H  v   x  `  w  w  x     y  ~  M   �     �M  �  �M    �M  �   �M  �  �M  �	  �M  �  ��   �    ��    ��  �  ��  �  ��   �  �  ��  �  ��  �  ��  m  �   �  	  �  2	  �  �  �  9  �  [  �Q   �  J  �Q  �  �Q  7  �Q  �  ��   �  I	  ��  $	  ��  �   ��   �  N  ��  p  ��   �  �  ��  :  ��  �  ��  d   ��  �  �   �    �  �  �  �	  �6   �  �  �6    �S   �  �  �S  �  �S  �  �S  +  �   �  �  �  �   �    �     �
  �  �  �    ��        ��  F  ��  �  �     �  �  �  �  �  3,   /  �  4,  �   8I   :  �  9I  l	  =f  E  N  >f  ^  ?f  L  @f  a  D�  P  B  E�  �	  F�    G�    H�  y  I�  �  	 �   [  �  	!�  �   W    ++CCUNGk   ++CCUNG�9  .f  �   q  ,     H   I�  I� � k  P     O� �?  �0   (  �     N   c  	� ��   �  �� �� u� l� �� V� �  Ç �/  	� �n   	M� �R   	$� �R   	�� �R   	Ŋ �u  
Ç ��   �   |  u   Ç �    |  �   �  �Ȅ �  #  |  �    �   �� �� R   H  N  %   n  N  n    I   &  ,g  ->   b� 1�  	<� 4%    	M� <N  	5� Dn   �� In  �  T n  %    Ԡ I�  �  T {  n  %    {  � kT    R    � uT    R    �� |�   *h  ��  -}  n  N  N  %     c  �  abi �>   std  t  int �   /  �   �  �  T WC  In  ,� I%     4  �  �  !h  �  j� �%   �� �n  �� �N  � �n   N  �  �  )  T {  WC  In  ,� I%     �   7  L  !h  L  �� �u   |  �  g  � kR      }  � uR    "#-  ���   �E  $� -n  � $�� .N  �$�� /N  �$j� 0%   �%� &`� 2n  L 'P� 3�  'X� 6n  &M� 8N  /L (�T  9�   �L)�  	� 77  *�  BL *�  aL  ))  �  9Z  +@  *7  �L  ,Q  Y�   ?w  *[  �L  ,Q  m�   B�  *[  �L  ,g  u�   F�  *q  VM  -�  ��8 M*�  �M .�  �*�  �M *�  �M *�  N ,�  ��   �  *�  5N *�  HN  /��   .�  S.�  �*�  gN .�  V.�  W    0   �   ��  � �� k  `     ̏ std  6  v  6�  x  K�  �  M6   x  Ob   m   8  6   	�  Qw  �   �   8   	�  R  �   �   8   
  T8  6  �   �   >   x  Z�   �   8   x  \�   �   8  D   x  _�     8  �   x  c  #  8  O   �  p�  U  ;  F  8  D   �  t�  U  ^  i  8  O   �  {y  �  8  [   n	 ~%  �  �  8  U   �  ��  b  �  �  >   �  �h  i  �  >    ;    :;   �  �J  � �  v�  w�  {�  ��  �  �   �5  �  ��  ��  ��  ��  �  �2  �S  �^  �o  ��  ��  ��  3�  �� �  �� ?�  Z    z �  z 9�  }    ��  �  ��  ��  �    v�   v� ��  �    ��   �� G  �    �� �� X.  		     ;   �  �  �  ;   ;   int �  �  �  (  _� 	Ԉ  �  	�  �  �  	��   �  	��   #  ��  
  	��  �  
�  �  �  o  �	  �  qW  
![    
"  �  s  N�  �  V�  .  <�  `  D[  �  W�  �  _
  �  e[  t   m[  a  u[    ~[  �  �[  3  �[  �  �[  H  �[  y  �[    �[  s  �[  T   �[  �  �[  F  �[  �  �[  �  �[    �[  V  �[  o  �  \	  2[  o  7[  �  <[  �  C[  �  [  !*  �  �  [   "rem [   +   h  !#@  �  �  $v   "rem %v   A  &�  #� �[  �  �   �  $#�  >�  �      ��   o  #�  H[         #�  Iv  5      #�  �6  ^  ^  ^  }  }  e   d  %k  &[    ^  ^   'div �  �  [  [   #    �$  �      (�   �  �  v  v   (�  .[  �     }   (�  \}         }       (3  >[  2       }   )�  S  6  }  }  e   *k� q[  +�  |o  �   #  W�  �     �   $  #  fv  �     �  [   #�  g�  �     �  [   #?  �[  �      �  =     =  ,��  !,p� %,�� ),�� --P  @m   ++CCUNG-}  Lm  ++CCUNG .abi ��  /T  6   I  �  0�  n  x  1h  x   Z  �  0�  �  �  1h  �   }  �  0�  �  �  1h  �   �  �  0�  �  �  1h  �   �    0
  �  	  1h  	   �    0"  	  '	  1h  '	   		  2�  ��#   �o	  3�  ��   "\	  4�  zN  5���  5��   2�  �#   ��	  3�  �   &�	  4�  �N  5��  53��   2  @�#   ��	  3�  M�   *�	  4�  �N  5J��  5c��   2  p�#   �8
  3	  }�   .%
  4	  �N  5z��  5���   6D  OD
     6�  PD
  61  QD
  6�  Wm
   '  6^  Xm
  6U  =�
   2  6�   >�
  6B  ?�
  6�  E�
   =  6B   F�
  6C  G�
  6e  H�
  68  I�
  6�  J�
  6

  X    H  6�  Y   6�
  Z   7�   `)  S  6�  f:   ^  6�  g:  6�  h:  6�  nc   i  6�	  oc  6�  pc  6H  v�   t  6`  w�  6w  x�  6   y�  6~  �     6   ��  6�  ��  6  ��  6�   ��  6�  ��  6�	  ��  6�  �   �  6  �  6  �  6�  �  6�  �O   �  6�  �O  6�  �O  6�  �O  6m  ��   �  6	  ��  62	  ��  6�  ��  69  ��  6[  ��   �  6J  ��  6�  ��  67  ��  6�  ��   �  6I	  ��  6$	  ��  6�   �#   �  6N  �#  6p  �@   �  6�  �@  6:  �@  6�  �@  6d   �@  6�  Ɂ   �  6  ʁ  6�  ˁ  6�	  Ѫ   �  6�  Ҫ  6  ��   �  6�  ��  6�  ��  6�  ��  6+  ��   �  6�  ��  6�   ��  6  �%     6�
  �%  6�  �%  6  �N     6   �N  6F  �N  6�  �w     6�  �w  6�  �w  6�  3�   1  6�  4�  6�   8�   <  6�  9�  6l	  =�  G  6N  >�  6^  ?�  6L  @�  6a  D  R  6B  E  6�	  F  6  G  6  H  6y  I  6�   \   ]  6�  !\  �  8   ++CCUNG8(  ++CCUNG9�  6  �  �   :�  6  6  T       ��  � 3� k  �     � �?  �0   (  �     �   �  	� ��   �  �� �� u� l� �� V� �  6� ��   	� ��   	�� �R   	.� ��  	�� ��  
6� ��   �  �    Ç ��  	� ��   	M� �R   	$� �R   	�� �R   	Ŋ ��  Ç �=  H  �  �   Ç �X  c  �  �   �  �Ȅ    w  �  �    �   �� � � �  I   �  �  �  �  0    I   �� �  �� !ˋ � W�   $  ,�  ->   �� I�    T �  %    �� |�   *�  � ��  �  I    �� ��  � �b  r      �   � +  �  �    �   � ��  �       �  �� $  �  �       �� +v� �  +  �    *  %   R   �  �  �  �      �  �� R   +  ;  U  *  %   �  �  �    �� J�� �  +  q  *  �  �  0    +   !�  �  "abi �>   #std  �  � �  U  x�� �  �  a  g    �   !�  $%int !�   !�   &�  &�   !+  !    �  &�  &+  !�  &�   'r  D  W  (h  W  (#  \     �  !�  &�  '�  {  �  (h  �  ):� x�   a  g  '  �  �  (h  �  )j� !%   )�� "�  )�� #�  )� $�   *  *�    T )WC  I�  ),� I%    'U    @  (h  �  +dst K�  )�� K�  )�T  L@   0  ,6  �� ��   �`  w  -D  � .��/� �   ,6  Ǣ ��!   ��  �  -D  � 06  ��   �  1D  �N 2�� 3���   4�  ��:  ��  �  5h  �  � 6j� ,%   �6� -R   �6�� .�  �6�� /�  �6�� 0�  �6� 1�  �6�T  2�  �0m  �.   4z  1{  �N 1�  O 7;�   0�  ��   9�  1�  ZO 1�  yO  8m  ��*   ?-{  U-�  �\7�       9�  ��  ��   ��  t  -�  � -�  �-�  �-�  �-�  �:� H  1�  �O 1�  �O 1�  �O 1�  �O 1�  P  8m  v�"   &1{  P 1�  :P 7��    9  �� ��Q   ��  �  -  � -  �-)  �-4  �:� �  14  YP 1)  xP 1  �P 1  �P  7���   �  ;  <�  1       =>mw  ww  �        �    ^�  �� T� k  ̔ (  �  �  int �  =D   �     �   �� %4� �   P  @�    ++CCUNG}  L�   ++CCUNG �  abi �K   	std  �   �� W�    
�   �  V   �D9   e    ++CCUNGy   ++CCUNG �   �  � �� k  `     ڕ �  (  _� �>   �  �  P   �  �  o  �	  pW   w   �  qW  !�   int   "�   �    #�   #  s  NE   �  VE   Fd ~   .  <~   `  D�   �  W~   �  _�   �  e�   t   m�   a  u�     ~�   �  ��   3  ��   �  ��   H  ��   y  ��     ��   s  ��   T   ȉ   �  Љ   F  ׉   �  ��   �  �     �   V  �   %   �  \	  2�   o  7�   �  <�   �  C�   �  �   E   	*  7  	�  	�    
rem 	�    +  	   	#@  g  	�  	$,    
rem 	%,    A  	&B  std    
v7  
wg  
{  
�  
�D  
�Y  
�n  
��  
��  
��  
�  
�  
�K  
�k  
��  
��  
��  
��  
��  
�  b�  c]  eh  f�  g�  h�  i�  j�  k�  l	  m-	  qG	  rl	  t�	  u�	  v�	  x�	  y�	  |	
  ~
  �0
  �E
  �_
  �q
  ��
  ��
  ��
  ��
  � �  H�  cÑ 9  �  �
    �  �� �   � 	��          �  	>2  2  9   �� ?  %   �  	H�   Y  9   �  	I,   n  9   �  	�   �  �  �  3   3   �   �  �  �   �  �  �   div 	7  �  �   �        	��  �  9   �  	 g    ,   ,    �  	.�     9  3    �  	\3   >  >  9  3    D    3  	>�   k  >  9  3    �  	�  �   3   3   �   k� 	q�   �  	|�  w      	W2  �  9  �   �    	f,   �  9  �  �    �  	g>     9  �  �    ?  	҉     9      W  D� ��  J  9  �  	     '� z�   �  abi �  	\  �   gX  �   X\  &�  X\  X,�  	$Z  .�    	\ /E   	� 1  	Z  23   	K]  3E   	�_  43   	\W  53   	�Z  63   	-_  8�   	VY  9�  $	`  :�  (	�Y  ;  ,	7_  <'  0	BY  =F  4	b\  >'  8	\  ?'  <	7Y  @'  @	 Z  AW  D	SX  BW  H	n4 Dl   L	`  F�  P	*5 G�  T u  �  �   3   �   �  �  u  �  �  3   �   �  �   �  �  j  �    �  j    �     �   '  �     �  F  9  9  �   -   W  �   L  �^  !j  Z  1z  z   �  aY  ��   �  z   \  C�   �  z   xZ  M�   �  z   `  ��   �  z   �^  r�   �  z   _X  ��   	  z  	   ]  �_  ��  -	  �  �   z   �\  �z  G	  9  9   4Z  �3   l	  �  3   3   z   7`  �z  �	  9  9  z   >]  	�   �	  z  ,   �    �Z  �   �	  z  �	   �	  ]  �Y   ,   �	  z   �Y  ��   �	  z   \  ��   �_  0�  
  �   �]  W0
  9   D[  T�   E
  9   �[  a�   _
  9  9   �\  )q
  z   Y@ ��
  z  �   �[     �
  z  �  �   3    �]  iz  D]  w�  �
  �   }W  ��   �
  �   z   !"r  !#  �  "�      #h     �
  $   �.  $�� ,S�  %"  �r  ��  &�j  �  '�� .W  �O(t 8�  �P )� �  *H�  <9  +�
  <� <�  ,  �P  )  �  '�� >�   �l(dem ?�  �P -[�&  -t�  -��;  -��  -��;  -��V   )H d  (exc R�  :Q &��A   H  (w T9  MQ -�  -*�;  -9�g   -���  -A��  -f��   -���  -x��  -���   -1�J  -��  -���  -F��  -Z�   -o��   �  �  .�  /D  O�   �   /�  P�  /1  Q�  /�  W�   �   /^  X�  /U  =   �   /�   >  /B  ?  /�  ED   �   /B   FD  /C  GD  /e  HD  /8  ID  /�  JD  /

  X�   �   /�  Y�  /�
  Z�  0�   `�  �   /�  f�     /�  g�  /�  h�  /�  n�     /�	  o�  /�  p�  /H  v     /`  w  /w  x  /   y  /~  R   #  /   �R  /�  �R  /  �R  /�   �R  /�  �R  /�	  �R  /�  ��   .  /  ��  /  ��  /�  ��  /�  ��   9  /�  ��  /�  ��  /�  ��  /m  �   D  /	  �  /2	  �  /�  �  /9  �  /[  �V   O  /J  �V  /�  �V  /7  �V  /�  ��   Z  /I	  ��  /$	  ��  /�   ��   e  /N  ��  /p  ��   p  /�  ��  /:  ��  /�  ��  /d   ��  /�  �   {  /  �  /�  �  /�	  �;   �  /�  �;  /  �X   �  /�  �X  /�  �X  /�  �X  /+  �   �  /�  �  /�   �  /  �   �  /�
  �  /�  �  /  ��   �  /   ��  /F  ��  /�  �   �  /�  �  /�  �  /�  31   �  /�  41  /�   8N   �  /�  9N  /l	  =k  �  /N  >k  /^  ?k  /L  @k  /a  D�  �  /B  E�  /�	  F�  /  G�  /  H�  /y  I�  /�   �     /�  !�  1F�  @z  3   �   2�� �� >   ;  �  3   3   z   �� ��   V  9  z     ;g  �    2�� �� �   �  �   z   3�  �   �  �    4�  4�  5f� 	�6>  Y  �     R   ��  �� *� k  �     w� (  �       A  P>�   �  AA   t  BR  +  F*  �  G5  �  J_  p  NB  p  YB    Ze  �  [e   �  \I  $w  ]  (4  a�  0 =  Ppx    s   �  xR  +  |*  �  }5  �  �_  p  �B  p  �B    �e  �  �e   �  �I  $w  �  (4  ��  0 �  ��  �  �_   �  �;   W  `  �  T   �  �  �  �   �  �_  �     	'� $A  
P  @6   ++CCUNG
}  L6  ++CCUNG�  X0   �  abi �3   + 0;  �  int (  5;  �  =_  �  B�  �  �   �  M  3  �  ]  K  	  �   �  Lf  �  W�  �  �  �  �   �  ^   Z  �  \T   �  ]�  V  b0  `  c0   std  A  � �� ZX  �� WX   %  R     G  ^  >   k  p  �  �  �  c `T   �   �  �  exc ��   �  �  ptr �   �  ��4   �0  p �  &0  vQ e  '_  �Q ��   %  de ,�   �  ��   .!�  �Q   "��    x  T  #�   ++CCUNG#�  ++CCUNG �    |�  �� b� k  �� (  �  �  int �  =D   �     �   �� � �   P  @�    ++CCUNG}  L�   ++CCUNG �  abi �K   	std  �   �� Z�    
�   �  V   �D9   e    ++CCUNGy   ++CCUNG �   !�  G�  � k  �     �� std  ~  v  6�  x  K�  �  M~   x  Ob   m   �  ~   	�  Qw  �   �   �   	�  R  �   �   �   
  T8  ~  �   �   �   x  Z�   �   �   x  \�   �   �  �   x  _�     �  �   x  c  #  �  �   �  p�  �  ;  F  �  �   �  t�  �  ^  i  �  �   �  {y  �  �  �   n	 ~%  �  �  �  �   �  ��  �  �  �  �   �  �h  �  �  �    ;    :;   �  ��  � �  �� Ux  n  n   �� X%  +  �   5� �  @  K  �  �   (�  a� �  �  g  �    z �  ��  ;   �  �  �  ;   ;   int �  �  �  �  �  �  s  +  �  �   h  �   #  �   �  �  !K  ��   �  $  "h  $  �  �  #�  � ��   �D  [  $�  � %��&� �   #�  � ��!   �v  �  $�  � '�  ��   �  (�  �Q )� *��   +�  �1  ~    Z   ��   � /� �V  @!     F� (  _� �7   �  �  8k  �{  k   ]�  k  \�   k  �D  !k  �3  "k  U>  #k  &�  $k  �  %k  �*  &k   ڡ  'q  $�U  (q  %TL  )q  &�I  *q  'Q  +q  (�C  ,q  )�J  -q  *1  .k  ,o(  /q  0�U  0q  1PL  1q  2�I  2q  3Q  3q  4�C  4q  5�J  5q  6 q  �  std ( .)  5>   6.)  7Z)  	Rk)  	U�)  	[�)  	\�)  
v�+  
w�+  
{�+  
��+  
�,  
�,  
�/,  
�y,  
��,  
��,  
��,  
��,  
�-  
�,-  
�M-  
�X-  
�i-  
��-  
��-  
��-  @�-  	%  0�=  �  �b  �q  Fe  �H)  
�3  �=  �  �3  �3   Z  eq �<-  �3  �  �3  �3   lt ��1  �3  �  �3  �3   ��  eF  H)  �  �3  �3     �K  �9      �3   �(  
!  �3  +  �3    �3   1  �A  �3  O  �3  �3     �5  �'  �3  s  �3  �3     �3  �A  �3  �  �3    Z   +  :  Z  �  �3   e  �C   �P  e  �  �3   �B  $6  �3  �  �3  �3   eof (�:  e  ?  ,N0  e  �3    _� �7   �?  �%   K  \�  .   �e  _  �4  c�3  �J  d4  ��  qs  y  4   ��  s�  �  4  4   W  y�  4  H)    ,  �J  p:  �B    ,   %  k   �B  �  �  @4  k  4   �B    @4  H)    �e  y?  [V  +    �G  !�   <  x,  �4  {K  �J  |W  �J  �/  `S  ��1  ~J  �:  �J  �?  �%  ��  �K  �   I  �  :!  �04   %H  �v  �   �3  2+  �G  7U)  t3  Bj4  �'  ��O  X4  V  ��N  �3    !  u4   3  �o+  �3  8  >  u4    �P  ��O  Q  W  R4    �M  ��P  j  p  R4    �,  �-  �  �  R4     �+  ��R  k  �  �  R4   3  �   k  �  �  R4  4  4   �/  !�B  R4  �      4    �O  �|6  	    R4  4   !(  ��6  (  3  R4  4   "�   �-  k  K  Q  R4   #�1  o�*  k  e  R4  4      "�A  $n%  k  �  �  F4   "�A  (�I  k  �  �  L4  k   ""A  ,�%  R4  �  �  F4   "�1  2E)  a  �  �  F4   "�/  6;&  a      F4   !�>  :�>  %  +  L4   "S  A:2    C  S  F4    O)   !�#  K�(  g  |  F4      O)   "9  S>$    �  �  F4       "-U  [�7  �3  �  �  F4  O)   $�5  d�-  �  k  O)     $	1  m�P  	  k  O)     $�3  v\-  '	  k    q   $nU  ��-  G	  k  a  a   $nU  �nG  g	  k  m  m   $nU  ��   �	  k  k  k   $nU  �IP  �	  k  O)  O)   �J  �rR  H)  �	       !�=  ��H  �	  �	  L4         !V  �)  
  	
  L4   %�'  �D*  X4  &�0  �*
  0
  L4   '�0  �@
  K
  L4  4   �0  �[
  f
  L4  ^4   �0  �v
  �
  L4  ^4       �0  ��
  �
  L4  ^4      4   �0  ��
  �
  L4  O)    4   �0  ��
  �
  L4  O)  4   �0  �
    L4    q  4   &�0  "0  ;  L4  H)   (�  *,Q  d4  T  _  L4  ^4   (�  2�G  d4  x  �  L4  O)   (�  =�%  d4  �  �  L4  q   (S� f�&  a  �  �  L4   (S� q�>  m  �  �  F4   )end y<  a  �    L4   )end �6;  m    #  F4   (I ��$  �  <  B  L4   (I ��7  y  [  a  F4   (��  �lC  �  z  �  L4   (��  �CM  y  �  �  F4   (r ��R    �  �  F4   (�K  �r5    �  �  F4   (�3  �j=    �  �  F4   *�� �    !  L4    q   *�� ��F  6  A  L4     (I  v    Z  `  F4   *�E  �|U  u  �  L4     *�1  -�  �  �  L4   (�� 5�?  �3  �  �  F4   (�:  D�6  U  �  �  F4     (�:  UW  I  �    L4     )at k
/  U    %  F4     )at ��7  I  =  H  L4     (�F  ��/  d4  a  l  L4  ^4   (�F  �k:  d4  �  �  L4  O)   (�F  ��H  d4  �  �  L4  q   (@  DA:  d4  �  �  L4  ^4   (@  U�1  d4  �    L4  ^4       (@  )�D  d4    /  L4  O)     (@  ��*  d4  H  S  L4  O)   (@  �6  d4  l  |  L4    q   *�G  -aN  �  �  L4  q   +�3  �b*  d4  �  �  L4  ^4   (�3  ^ 2  d4  �  �  L4  ^4       (�3  �=  d4      L4  O)     (�3  z�T  d4  /  :  L4  O)   (�3  � @  d4  S  c  L4    q   *� ��E  x  �  L4  a    q   (� �\+  d4  �  �  L4    ^4   (� �u>  d4  �  �  L4    ^4       (� g|=  d4      L4    O)     (� "�@  d4  0  @  L4    O)   (� 9k<  d4  Y  n  L4      q   (� K�'  a  �  �  L4  a  q   (bL  d�R  d4  �  �  L4       (bL  t�2  a  �  �  L4  a   (bL  �L&  a  �    L4  a  a   (�%  �9F  d4  &  ;  L4      ^4   (�%  �|<  d4  T  s  L4      ^4       (�%  ��T  d4  �  �  L4      O)     (�%  ��A  d4  �  �  L4      O)   (�%  b>  d4  �    L4        q   (�%  3%  d4     5  L4  a  a  ^4   (�%  'V7  d4  N  h  L4  a  a  O)     (�%  <�+  d4  �  �  L4  a  a  O)   (�%  Q'S  d4  �  �  L4  a  a    q   (�%  vj.  d4  �  �  L4  a  a  k  k   (�%  ��9  d4    /  L4  a  a  O)  O)   (�%  �C  d4  H  b  L4  a  a  a  a   (�%  �>/  d4  {  �  L4  a  a  m  m   "�?  ��&  d4  �  �  L4        q   "�1  �O  d4  �  �  L4      O)     ,)  �z-  k      q  4   ,+E  �3J  k  @    q  4   (�5  ��)    Y  n  F4  k       *n	 @D  �  �  L4  d4   (W�  �6  O)  �  �  F4   (�A  %�A  O)  �  �  F4   (��  ,Z5  =  �  �  F4   (�(  �;        F4  O)       (�(  I�%    2  B  F4  ^4     (�(  X�5    [  k  F4  O)     (�(  �^     �  �  F4  q     (�(  v�S    �  �  F4  ^4     (�(  	K    �  �  F4  O)       (�(  �o?        F4  O)     (�(  J5    -  =  F4  q     (NW  ��Q    V  f  F4  ^4     (NW  /�I      �  F4  O)       (NW  ��,    �  �  F4  O)     (NW  ��;    �  �  F4  q     (�S  ��I    �    F4  ^4     (�S  >T?    (  =  F4  O)       (�S  05    V  f  F4  O)     (�S  $S:      �  F4  q     (�>  2hL    �  �  F4  ^4     (�>  SUB    �  �  F4  O)       (�>  Q�2    �    F4  O)     (�>  _�K    (  8  F4  q     (�4  qT    Q  a  F4  ^4     (�4  j�K    z  �  F4  O)       (�4  ��5    �  �  F4  O)     (�4  N.    �  �  F4  q     (U+  �)  �  �  
  F4       (��  �!1  H)  #  .  F4  ^4   (��  ��T  H)  G  \  F4      ^4   (��  ��O  H)  u  �  F4      ^4       (��  �;.  H)  �  �  F4  O)   (��  ��B  H)  �  �  F4      O)   (��  ��,  H)  �    F4      O)     �  -!T  q  .�E  N  .�F  ,   /�&  /�7  �  �o  >#  �| CH)  0Q  bn   U  0�F cn  0�R  dn  03  en  0�  fn  0�K  gn  0�@  hn   1all in  ?2�� �   :!  �04   NF  ��4  �E  �  p0  ��4  �%  ��-  3S  ��4  3�R  ��4  33  ��4  3�$  ��4  3�K  ��4  3�@  ��4  3�@  ��4  !�4  �Z  �  �  {4   !�=  y)  �  �  {4   �� �  �  {4  �4     �� �  �  {4  O)     �� �     {4     N      {4  H)   �� +  6  {4  �4   !�  �U  J  U  {4  �4   "�&  �.  �3  m  s  {4   !�F  &�;  �  �  {4  �4  U   !�9  )�Q  �  �  {4  �4  �4   !WR  ,`2  �  �  {4  �4  �4   !�S  /=  �    {4  �4  �4   !e  7,    '  {4  �4     �� 3@  K  -�R  F$  {4  �:   � 3d  o  -�R  \$  {4  5;   � 3�  �  -�R  �$  {4  �;   � 3�  �  -�R  	%  {4  �;   �� 3�  �  -�R  M%  {4  &<   � 3�  �  -�R  �%  {4  �<   �� 3  #  -�R  �%  {4  �<   � 3<  G  -�R  D&  {4  �<   +� 3`  k  -�R  �&  {4  =   ƪ 3�  �  -�R   '  {4  w=   E� 3�  �  -�R  D'  {4  �=   &� 3�  �  -�R  c'  {4  >   �� 3�  �  -�R  �'  {4  b>   4�� 3   -�R  �'  {4  �>    �$  {4   3OD  {4  3gP  {4  3�F  $�4  5< �   6< rg   r   �9     7�m  �~�  ")  7��  ���  O)   8id �&!  �U  �   3�I  �04  !�  �<?  �   �   �4  �4   9id ��   �   �4  �4   :id �!  
!  �4   ;4H  ��(    !  �4    �o  u6!  <!  �4   �o  ~L!  W!  �4  �4   '�o  �g!  r!  �4  O)   �o  ��!  �!  �4  �4  O)  U   �o  ��!  �!  �4  �4  �4  U   5  ��!  �!  �4  H)   +�  ��*  �4  �!  �!  �4  �4   +H�  ��N  #  "  "  �4   +U  �9  �3  0"  ;"  �4  �4   +2  �t*  �3  S"  ^"  �4  �4   <jP  �D  I  y"  �4   7RD  �Q  �4  =�o  7�"  �"  �4  {4   >�K  :�N  >�A  =�5  �K  @I  U  �"  U   !�,  CH<  �"   #  �4  �4  �4  U   �   M   �   I  � >�  <�4  =�4  >5  @�5  A�5  B�5  C�5  D�5  E6  F/6  GD6  HY6  ks  4�#  ?ks  �#  �:    @�  H$  ASv  L�#  �O  L}6    �  N�#  �#  ��  YO)  <Fv  ^��  �#  �#  q  q  q   ?�  $  �:    ד  �F$  ��  �!  � �k  �4  ��3  -{�  k   5�+  \$  Bid ��    5(�  r$  Bid a�    C0T  �$  ��  :�$  �$  h;     -!T  q   5�N  	%  6��  ��$  �$  �;  QA     D��  rr$  Bid >�   -!T  q  E��  E��  �$  �;  ")    5�p  M%  6mF �#%  .%  �;     Bid ��   -!T  q  .�  )   5"(  �%  6H �g%  r%  &<     Bid �	�   -!T  q  .QJ  )   5_}  �%  63  c�%  �%  �<     Bid ��   -!T  q   5��  D&  6�q  ��%  �%  �<  �A     D��  �v(  Bid �   -!T  q  F�  �3   E�q  ��  3&  �<  ")  O)    5�  �&  6�q  �^&  n&  �<  NB     D��  ��(  Bid �   -!T  q  F�  �3  E�q  Y�  �&  �<  ")  O)    5��   '  6��  p�&  �&  =     Bid ��   -!T  q  .�  )   5�  D'  60�  '  %'  w=     Bid |�   -!T  q  .QJ  )   5��  c'  Bid B�   -!T  q   5C�  �'  6��  �}'  �'  >     Bid ��   -!T  q  .�  )   5|  �'  6�p  ��'  �'  b>     Bid '�   -!T  q  .QJ  )   5l�  
(  Bid H�   -!T  q   G&� �	�3  @(  -!T  q  -�E  N  -�F  ,  ^4  O)   G�� 
�3  v(  -!T  q  -�E  N  -�F  ,  ^4  O)   C
�  �(  ҽ  z�(  �(  �A     -!T  q  F�  �3    C��  �(  ҽ  z�(  �(  B     -!T  q  F�  �3   C�  )  H�  z�(  	)  �B     -!T  q   #  /��  /;G  W�  1�Y   I)%  Kk  H)  H)  O)   Jint U)  q  KGT  Pe)  >   I��  EH)  �)  O)  O)   I��  Uk  �)  H)   I��  Ok  �)  k  O)   I��  F,   �)  k  O)  ,    �  �)  �  �  o  �	  �  qW  !H)    "*  �  #  Ls  N�)  �  V�)  .  <*  `  DH)  �  W*  �  _*  �  eH)  t   mH)  a  uH)    ~H)  �  �H)  3  �H)  �  �H)  H  �H)  y  �H)    �H)  s  �H)  T   �H)  �  �H)  F  �H)  �  �H)  �  �H)    �H)  V  �H)  �  \	  2H)  o  7H)  �  <H)  �  CH)  �  H)  M*  �+  �  H)   Nrem H)   +   m+  M#@  �+  �  $%    Nrem %%    A  &�+  I� �H)  �+  �+   �+  OI�  >�+  �+  O)   �� I�  HH)  ,  O)   I�  I%   /,  O)   I�  �%*  X,  X,  X,  ,   ,   _,   ^,  Pe,  QH)  y,  X,  X,   Rdiv �+  �,  H)  H)   I    �k  �,  O)   G�   �+  �,  %   %    G�  .H)  �,  O)  ,    G�  \,   �,  �,  O)  ,    -    G3  >H)  ,-  �,  O)  ,    S�  M-  %*  ,   ,   _,   Kk� qH)  T�  |i-  �)   I  W�+  �-  O)  �-   k  I  f%   �-  O)  �-  H)   I�  g7   �-  O)  �-  H)   I?  �H)  �-  O)   UpO qO !�-  V$   #E�3  	�  $ ,   -!  K   :�/  �e   =  �  ?k  "   @O)  �4   A�3  �J   B4  �A   Og.  m.  4   �A   Q}.  �.  4  4   �A   V�.  �.  4  H)   +�
  Y51  '.  �.  �.  4  ?.   +�
  ]�R  3.  �.  �.  4  K.   +�  c?  '.  /  /  4  .  X,   W_  m.   %/  5/  4  '.  .   +�3   q89  .  M/  S/  4   W.E   ��3  g/  w/  4  '.  4   W�(   ��(  �/  �/  4  '.   X_Tp q   .  @ZD  !��1  YF�  !�k   D��  !�$  D�4  !�1$  D� !�&$  &��  !��/  �/  �6   6��  !�0  0  �6  �6   (*  !��}  �/  30  90  �6   (Ư  !�?s  �/  R0  X0  �6   (�F  !�Ϭ  �6  q0  w0  �6   (�F  !��  �/  �0  �0  �6  H)   (a�  !�
�  �6  �0  �0  �6   (a�  ! ��  �/  �0  �0  �6  H)   (�:  !,�  �/  �0  1  �6  �/   (�F  !		n  �6  1  &1  �6  �/   ((*  !��  �/  ?1  J1  �6  �/   ( I  !h�  �6  c1  n1  �6  �/   (�O  !7k  �/  �1  �1  �6  �/   (WC  !]�  �6  �1  �1  �6   -{�  k  -�  �   /8E  �/  Z*; "1�1  [�8  [�; [N;  �; "v�2  �= "|%4   H�; "2  2  �6  �6   �  "��= �6  62  A2  �6  �6   �; "�Q2  W2  �6   W\ "��: k2  q2  �6   Wf "��8 �2  �2  �6   \�9 "��: �6  �2  �6    �1  (8 "�>3  r< "��1  �9 "��6   H(8 "��2  �2  �6  �6   �  "�< �6   3  3  �6  �6   '(8 "�3  &3  �6  �6   '8 "�23  �6  H)    �2  ]U  A04  ]3  �8  H)   ^��  Is3  �8  H)   ]9+  N04  �3  �8  H)   ^��  \�3  �8  H)   _�= "5�3   �1   �� �� V2*  7�3  `8G   aZ  a�  �  �  Z  a�  aq  aU)  .  a�/  �/  ,  a�  ��  $!H)  �  % H)  H)  �  D  �  �  a�  aD  a�  b7   u4  c   �  �4  �4  O)  I  a#  #  �   a #   #  �4  #  b�4  �4  c b�4  �4  c �4  �4  a
#  
#  �l  &%   j�  &#%   dtm ,&,�5  ,g  &.H)   �  &/H)  �  &0H)  ��  &1H)  ��  &2H)  ��  &3H)  ��  &4H)  �  &5H)  d�  &6H)   ��  &7%   $~�  &8O)  ( K\�  &>�4  Iѯ  &H�+  �5  �4  �4   I��  &M�4  �5  �5   5  I�  &C�4  �5  �5   �4  I#�  &ak  6  6   
6  5  I�� &fk  $6  $6   *6  �4  I��  &W�5  D6  $6   I[v  &\�5  Y6  $6   I��  &R,   }6  k  ,   O)  6   bq  �6  e/+   �/  a�6  k  �1  a�/  �1  a�2  a�1  %4  �6  a�2  �2  a>3  a�2  f�8  `(x  g�� "�6  � *ZW  h-� ,�6  � .}6  h8 07  hn� 4�W  h� 8�W  h� <�W  h;� @�W  � B�W  h� DN7  ڮ FX  h߮ Hd7  � JX  h� Lz7  �� N:X  hĭ P�7  � R:X  h� T�7  � VX  h!� X�7  {� ZX  hX� \�7  hJ� ]�7  î _:X  hȮ a�7  n� c:X  hs� e	8  �� gZW  h�� i8  �� k:X  h�� m58  � o:X  h$� qK8  �� s�X  h�� ua8  �� ��X  h�� �w8  l� ��X  hذ ��8  hg� ��8  � �"Y  h� ��8   ` �6  04  iC3   9  jXF  A�8  j\;  AH)  kl�T  C04    i]3  !9  jXF  I�8  j\;  IH)   mv  /9  99  nh  99   F4  i�  V9  ko__p �%*    is3  w9  jXF  N�8  j\;  NH)   m�  �9  �9  nh  �9  p__a �9   R4  4  q�  '�%*  �9    p__p '�%*   q�  '�%*  �9    p__p '�%*   r�  '��9  %*  %*   M   mV   :  ':  nh  ':  s4&  r   �9  i�3  M:  jXF  \�8  j\;  \H)   mA2  [:  e:  nh  e:   �6  i�6  �:  kl�� $�1    mW2  �:  �:  nh  e:   mq2  �:  �:  nh  e:   �#  t�#  H�:  �:  nh  �:   �:  t#  u�#  4�:  �:  nh  �:   �:  F$  m'  ;  0;  -�R  F$  nh  0;  sf� 3�:   {4  \$  mK  R;  h;  -�R  \$  nh  0;  sf� 35;   r$  m{$  |;  �;  nh  �;  s4&  :   h;  �$  mo  �;  �;  -�R  �$  nh  0;  sf� 3�;   	%  m%  �;  �;  nh  �;  s4&  �   �;  m�  <  &<  -�R  	%  nh  0;  sf� 3�;   M%  mV%  :<  P<  nh  P<  s4&  �   &<  m�  l<  �<  -�R  M%  nh  0;  sf� 3&<   �%  m�  �<  �<  -�R  �%  nh  0;  sf� 3�<   �%  m�  �<  �<  -�R  �%  nh  0;  sf� 3�<   D&  m#  =  =  -�R  D&  nh  0;  sf� 3�<   �&  m�&  /=  E=  nh  E=  s4&  p   =  mG  a=  w=  -�R  �&  nh  0;  sf� 3=    '  m	'  �=  �=  nh  �=  s4&     w=  mk  �=  �=  -�R   '  nh  0;  sf� 3w=   D'  m�  �=  >  -�R  D'  nh  0;  sf� 3�=   c'  ml'  >  0>  nh  0>  s4&  �   >  m�  L>  b>  -�R  c'  nh  0;  sf� 3>   �'  m�'  v>  �>  nh  �>  s4&  �   b>  m�  �>  �>  -�R  �'  nh  0;  sf� 3b>   �'  m�  �>  �>  -�R  �'  nh  0;  sf� 3�>   v�"  v�"  mq  ?  ?  nh  0;   m3  )?  >?  nh  >?  jF�  "�C?   �6  �6  m&3  V?  i?  nh  >?  n#  ;4   i
(  �?  -!T  q  -�E  N  -�F  ,  s\C  �	�?  s?)  �	O)   ^4  m�.  �?  �?  nh  �?  n#  ;4   4  m�  �?  �?  nh  �?  n#  ;4   4  mm.  @  @  nh  �?  @   4  my  (@  =@  nh  �?  p__a s=@   4  m�  P@  Z@  nh  99   m�  h@  r@  nh  99   t�  �@  �@  nh  �@  n#  ;4   @4  i@(  �@  -!T  q  -�E  N  -�F  ,  s\C  
�@  s?)  
O)   ^4  m�  �@  �@  nh  99   m  A  A  nh  A  n#  ;4   L4  wj:   �(   �QA  x#�!   yu:  z-��Y  zA��Y    �$  m�$  eA  �A  nh  �A  s��  �QA  s4&  �   �;  m�%  �A  �A  nh  �A  s4&  c   �<  v(  m(  �A  �A  nh  �A  s4&  z   �A  �%  m�%  �A  B  nh  B  s��  ��A  s4&  �   �<  �(  m�(  3B  IB  nh  IB  s4&  z   B  n&  mM&  bB  �B  nh  �B  s��  �NB  s4&  �   �<  �(  m�(  �B  �B  nh  �B  j4&  z   �B  t�  u �B  xC  nh  0;  s4&  v  k{�� �r$  |Ԯ ��B  �B  {�� �v(  {�� ��(  |�� � C  �B  |� �2C  C  {� ��(  |� �PC  8C  }hC  ~__i |   k~__j �     �B  P� P��  ��C  �K  ��B  � ��B  ��� �K  ��B  �Q �C  R �&C  RR �DC  zR ���   �C  �[C  �R  ���!   D  yiC   �;  	�   �7D  �#;  �R �;  �R z��   �;;  *�   �jD  �[;  US �R;  }S z:��   �WA  <�� ��D  �zA  T �nA  �Q �eA  $T �:  ��
   ��D  �:  T �:  $T  z���$  ��� �n;  C�l   �'E  ��;  LT �|;  lT �:  C�
   ?�:  LT �:  lT   ��;  ��   �ZE  ��;  �T ��;  �T z���   ��;  ��   ��E  ��;  <U ��;  hU �:  ��
   ��:  <U �:  hU   ��;  ��   ��E  �<  �U �<  �U z��   �,<  �   �-F  �C<  HV �:<  tV �:  �
   ��:  HV �:  tV   �U<  #�   �`F  �u<  �V �l<  �V z3��   ��A  6� ��F  ��A  TW ��A  �W �:  6�
   d�F  �:  TW �:  �W  zO�r   ��� ��<  O�( ��F  ��<  �W ��<  �W zg��   ��A  j�@ �FG  ��A  IX ��A  uX �:  j�
   ��:  IX �:  uX   ��A  ~�X ��G  �B  �X �B  R ��A  �X �:  5�
   ��G  �:  �X �:  �X  zX�"&  �� ��<  [�   ��G  ��<  Y ��<  9Y zk��   �%B  n�x �6H  �<B  {Y �3B  �Y �:  n�
   ��:  {Y �:  �Y   �TB  ��� ��H  �wB  �Y �kB  RR �bB  �Y �:  9�
   ��H  �:  �Y �:  �Y  z\��&  ��� ��<  _�   ��H  �=  Z �=  #Z zo��   �!=  r�   �&I  �8=  NZ �/=  bZ �:  r�
   p�:  NZ �:  bZ   �J=  ��   �YI  �j=  zZ �a=  �Z z���   �}=  ��   ��I  ��=  �Z ��=  �Z �:  ��
   �:  �Z �:  �Z   ��=  ��   ��I  ��=  �Z ��=  [ z���   ��B  ��� �+J  ��B  ,[ ��B  @[ �:  ��
   ��:  ,[ �:  @[   ��=  ��   �^J  ��=  X[ ��=  p[ z���   �>  ��   ��J  �#>  �[ �>  �[ �:  ��
   ��:  �[ �:  �[   �5>  ��   ��J  �U>  �[ �L>  �[ z���   �h>  ��   �1K  �>  
\ �v>  \ �:  ��
   ��:  
\ �:  \   ��>  �   �dK  ��>  6\ ��>  N\ z#��   ��>  4�   ��K  ��>  y\ ��>  �\ zD��   z���   ���'�����1�zS�
!  zi�
!  z�
!  z��
!   z���Y  z%�Z   ��>  �5  0�'   �L  z?�xC   w�>  `�'   �AL  ��>  c�    zo�xC    ��>  �N  ��   �dL  ���L   u&!  � tL  �L  nh  �L  kl�_ �2    �4  dL  � ��g   ��L  �M  �tL  � ��>  ��� ��L  z�L   �� zM  y~L  �j:  ��� �M  ���	   	M  yu:   z��A   �?  ��   �?  �\ �,:  ��   ��A:  �\ �6:  �\ � 9  ��   d�9  �\ �
9  �\     �?   �   ߅?  �\ �,:   �   ��A:  �\ �6:  �\ � 9   �   d�9  �\ �
9  �\     �y"    �<   �N  ��>  #�  N  zU�L   �:� �^"  �`�  ��Q  ��< �Q  ��(  �Q  �'U  �{4  
] ��>  i�H  �{N  z5�L   �h  �Q  l�_ �2  �� �)  �\�j:  z��  ��N  �z�	   �N  yu:   z��A   �?  ��   �;O  �?  3] �,:  ��   ��A:  F] �6:  3] � 9  ��   d�9  F] �
9  3]    ��@  ��   �O  ��@  r] ��@  �] �i?  ��   
��?  r] ��?  �] z���    ��@  ���  �P  �A  ^ �Z@  ���  #�O  �h@  ^ �!9  ���  -�/9  ^   �w9  ���  #��9  '^ ��9  I^ x�"   ��9  g^ ��9  �^ �V9  �! ��P  �k9  �^ �`9  �^ ��8  �! V��8  �^ ��8  �^ �! ��8  �^    z(�     ��@  :�7   �Q  �A  ud��Z@  :�   #�P  �h@  ud��!9  :�   -�/9  ud�  �w9  B�/   #��9  uc���9  �^ xS�   ��9  _ ��9  <_ �V9  S�(! ��Q  �k9  �`9  O_ ��8  S�(! V��8  ��8  O_ �(! ��8  S   zl�     z���!  z��.)   ��� zS��Y   �4  �D  O�Q   '*  ��  P�Q  �1  Q�Q  ��  W�Q   2*  �^  X�Q  �U  =R   =*  ��   >R  �B  ?R  ��  EFR   H*  �B   FFR  �C  GFR  �e  HFR  �8  IFR  ��  JFR  �

  X�R   S*  ��  Y�R  ��
  Z�R  ��   `�R  ^*  ��  f�R   i*  ��  g�R  ��  h�R  ��  nS   t*  ��	  oS  ��  pS  �H  v/S   *  �`  w/S  �w  x/S  �   y/S  �~  hS   �*  �   �hS  ��  �hS  �  �hS  ��   �hS  ��  �hS  ��	  �hS  ��  ��S   �*  �  ��S  �  ��S  ��  ��S  ��  �T   �*  ��  �T  ��  �T  ��  �T  �m  �:T   �*  �	  �:T  �2	  �:T  ��  �:T  �9  �:T  �[  ��T   �*  �J  ��T  ��  ��T  �7  ��T  ��  ��T   �*  �I	  ��T  �$	  ��T  ��   ��T   �*  �N  ��T  �p  �U   �*  ��  �U  �:  �U  ��  �U  �d   �U  ��  �JU   �*  �  �JU  ��  �JU  ��	  �vU   �*  ��  �vU  �  ؕU   �*  ��  ٕU  ��  ڕU  ��  ەU  �+  ��U   +  ��  ��U  ��   ��U  �  ��U   +  ��
  ��U  ��  ��U  �  �&V   +  �   �&V  �F  �&V  ��  �RV   $+  ��  �RV  ��  �RV  ��  3~V   6+  ��  4~V  ��   8�V   A+  ��  9�V  �l	  =�V  L+  �N  >�V  �^  ?�V  �L  @�V  �a  D�V  W+  �B  E�V  ��	  F�V  �  G�V  �  H�V  �y  I�V  ��   HW   b+  ��  !HW  bq  jW  e/+   �7  �U�7  �Ubq  �W  e/+  e/+   �"7  �Ubq  �W  e/+  e/+   �-7  �Ubq  �W  e/+  e/+   �87  `U�C7   Ubq  X  �/+   �Y7   Sbq  "X  e/+   �o7  �R��7  �Rbq  JX  e/+   ��7  �R��7  �R��7  �R��7  �R��7  �R��7  �R�8  �R�*8  �R�@8  �R�V8  xRbq  �X  e/+   �l8  hRbq  �X  e/+  g ��8   Rbq  
Y  e/+  C ��8  �Q��8   Qbq  2Y  e/+  � ��8   P��3   �  w� l	�)  (�� \	�5  6�� T	�A  @� D	�M  Nέ 0	�Y  ^�� (	�e  hf� 	�e= H)  �Y  �Y   *  �Y< �Y  �Y   H)  �>  Y  Z  %*   �  %*    ),   @�  �� C� �V  �!     �� (  �  �  �  E   �  �  o  �	  �  qW  !s   int   "�   �  #  .  <h   `  Ds   �  Wh   �  _z   �  es   t   ms   a  us     ~s   �  �s   3  �s   �  �s   H  �s   y  �s     �s   s  �s   T   �s   �  �s   F  �s   �  �s   �  �s     �s   V  �s   3   �  s  N:   �  V:   \	  2s   o  7s   �  <s   �  Cs   �  s   �  �  3   		pO qO 	!�  
std  �  @�  %  0�=  
��  �b  
�3   Fe  
�s   �3  
�=  [  �   �    +  eq 
�<-  �   }  �   �    lt 
��1  �   �  �   �    ��  
eF  s   �  �   �   �   �K  
�9  �  �  �    �(  

!  �   �  �   �  �    1  
�A  �      �   �   �   �5  
�'  �   D  �   �   �   �3  
�A  �   h  �   �  +   +  
:  +  �  �    6  �C  
 �P  6  �  �    �B  
$6  �   �  �   �    eof 
(�:  6  ?  
,N0  6  �     _� �,   5�   6�!  7"  �?  �%   K  \�  �   �e  _�  �4  c("  �J  d."  ��  qY  _  F"   ��  so  z  F"  L"   W  y�  F"  s       �J  p   �B  �     %  �   �B  �  �  ^"  �  L"   �B  �  ^"  s     �e  y%  [V    �  �G  !�   <  x  �4  {1  �J  |=  �J  =   `S  �B   ~J  �   �J  �%  �%  ��   �K  ��    I  ��   :!  �"   %H  �\  w   !�3  2  !�G  7�  !t3  B�"  "�'  ��O  v"  #V  ��N  �       �"   #3  �o+  �     $  �"   $�P  ��O  7  =  p"   $�M  ��P  P  V  p"   $�,  �-  i  t  p"  �   #�+  ��R  �  �  �  p"   #3  �   �  �  �  p"  L"  L"   �/  !�B  p"  �  �  �  L"   $�O  �|6  �  �  p"  L"   %(  ��6      p"  L"   &�   �-  �  1  7  p"   '�1  o�*  �  K  p"  L"  �    &�A  $n%  �  t  z  d"   &�A  (�I  �  �  �  j"  �   &"A  ,�%  p"  �  �  d"   &�1  2E)  G  �  �  d"   &�/  6;&  G  �  �  d"   %�>  :�>      j"   &S  A:2  �  )  9  d"  �  �   %�#  K�(  M  b  d"  �  �  �   &9  S>$  �  z  �  d"  �  �   &-U  [�7  �   �  �  d"  �   (�5  d�-  �  �  �  �   (	1  m�P  �  �  �  �   (�3  v\-  	  �  �  3    (nU  ��-  -	  �  G  G   (nU  �nG  M	  �  S  S   (nU  ��   m	  �  �  �   (nU  �IP  �	  �  �  �   �J  �rR  s   �	  �  �   %�=  ��H  �	  �	  j"  �  �  �   %V  �)  �	  �	  j"   )�'  �D*  v"  *�0  �
  
  j"   +�0  �&
  1
  j"  L"   �0  �A
  L
  j"  |"   �0  �\
  q
  j"  |"  �  �   �0  ��
  �
  j"  |"  �  �  L"   �0  ��
  �
  j"  �  �  L"   �0  ��
  �
  j"  �  L"   �0  ��
    j"  �  3   L"   *�0  "  !  j"  s    ,�  *,Q  �"  :  E  j"  |"   ,�  2�G  �"  ^  i  j"  �   ,�  =�%  �"  �  �  j"  3    ,S� f�&  G  �  �  j"   ,S� q�>  S  �  �  d"   -end y<  G  �  �  j"   -end �6;  S    	  d"   ,I ��$  k  "  (  j"   ,I ��7  _  A  G  d"   ,��  �lC  k  `  f  j"   ,��  �CM  _    �  d"   ,r ��R  �  �  �  d"   ,�K  �r5  �  �  �  d"   ,�3  �j=  �  �  �  d"   .�� �  �    j"  �  3    .�� ��F    '  j"  �   ,I  v  �  @  F  d"   .�E  �|U  [  f  j"  �   .�1  -�  {  �  j"   ,�� 5�?  �   �  �  d"   ,�:  D�6  ;  �  �  d"  �   ,�:  UW  /  �  �  j"  �   -at k
/  ;       d"  �   -at ��7  /  #  .  j"  �   ,�F  ��/  �"  G  R  j"  |"   ,�F  �k:  �"  k  v  j"  �   ,�F  ��H  �"  �  �  j"  3    ,@  DA:  �"  �  �  j"  |"   ,@  U�1  �"  �  �  j"  |"  �  �   ,@  )�D  �"      j"  �  �   ,@  ��*  �"  .  9  j"  �   ,@  �6  �"  R  b  j"  �  3    .�G  -aN  w  �  j"  3    /�3  �b*  �"  �  �  j"  |"   ,�3  ^ 2  �"  �  �  j"  |"  �  �   ,�3  �=  �"  �  �  j"  �  �   ,�3  z�T  �"       j"  �   ,�3  � @  �"  9  I  j"  �  3    .� ��E  ^  s  j"  G  �  3    ,� �\+  �"  �  �  j"  �  |"   ,� �u>  �"  �  �  j"  �  |"  �  �   ,� g|=  �"  �  �  j"  �  �  �   ,� "�@  �"    &  j"  �  �   ,� 9k<  �"  ?  T  j"  �  �  3    ,� K�'  G  m  }  j"  G  3    ,bL  d�R  �"  �  �  j"  �  �   ,bL  t�2  G  �  �  j"  G   ,bL  �L&  G  �  �  j"  G  G   ,�%  �9F  �"    !  j"  �  �  |"   ,�%  �|<  �"  :  Y  j"  �  �  |"  �  �   ,�%  ��T  �"  r  �  j"  �  �  �  �   ,�%  ��A  �"  �  �  j"  �  �  �   ,�%  b>  �"  �  �  j"  �  �  �  3    ,�%  3%  �"      j"  G  G  |"   ,�%  'V7  �"  4  N  j"  G  G  �  �   ,�%  <�+  �"  g  |  j"  G  G  �   ,�%  Q'S  �"  �  �  j"  G  G  �  3    ,�%  vj.  �"  �  �  j"  G  G  �  �   ,�%  ��9  �"  �    j"  G  G  �  �   ,�%  �C  �"  .  H  j"  G  G  G  G   ,�%  �>/  �"  a  {  j"  G  G  S  S   &�?  ��&  �"  �  �  j"  �  �  �  3    &�1  �O  �"  �  �  j"  �  �  �  �   ,)  �z-  �    �  3   L"   0+E  �3J  �  &  �  3   L"   ,�5  ��)  �  ?  T  d"  �  �  �   .n	 @D  i  t  j"  �"   ,W�  �6  �  �  �  d"   ,�A  %�A  �  �  �  d"   ,��  ,Z5  #  �  �  d"   ,�(  �;  �  �  �  d"  �  �  �   ,�(  I�%  �    (  d"  |"  �   ,�(  X�5  �  A  Q  d"  �  �   ,�(  �^   �  j  z  d"  3   �   ,�(  v�S  �  �  �  d"  |"  �   ,�(  	K  �  �  �  d"  �  �  �   ,�(  �o?  �  �  �  d"  �  �   ,�(  J5  �    #  d"  3   �   ,NW  ��Q  �  <  L  d"  |"  �   ,NW  /�I  �  e  z  d"  �  �  �   ,NW  ��,  �  �  �  d"  �  �   ,NW  ��;  �  �  �  d"  3   �   ,�S  ��I  �  �  �  d"  |"  �   ,�S  >T?  �    #  d"  �  �  �   ,�S  05  �  <  L  d"  �  �   ,�S  $S:  �  e  u  d"  3   �   ,�>  2hL  �  �  �  d"  |"  �   ,�>  SUB  �  �  �  d"  �  �  �   ,�>  Q�2  �  �  �  d"  �  �   ,�>  _�K  �      d"  3   �   ,�4  qT  �  7  G  d"  |"  �   ,�4  j�K  �  `  u  d"  �  �  �   ,�4  ��5  �  �  �  d"  �  �   ,�4  N.  �  �  �  d"  3   �   ,U+  �)  �  �  �  d"  �  �   ,��  �!1  s   	    d"  |"   ,��  ��T  s   -  B  d"  �  �  |"   ,��  ��O  s   [  z  d"  �  �  |"  �  �   ,��  �;.  s   �  �  d"  �   ,��  ��B  s   �  �  d"  �  �  �   ,��  ��,  s   �  �  d"  �  �  �  �   �  1!T  3   2�E    2�F     3�&  3�7  �  � >�  4W  3�  5�4  5�$  5q-  5c=  5o'  5�5   5�%  � 5�8  �5X)  �5�%  �5�  �5aO  �5Y=  � 5P  �� 5�C  ��5wS  �5�O  � 5�?  �5�5  �� 4
$ g  5)W  5�   5�U  5�A  5�8  5�P   5EH  �� 4�4  �/  5O   5�7  5(  5�Q  5G  �� 6b4 e  7�� �e  �  e    K� �/  8�� j  u  �"  �"   +�� #�  �  �"  �"   9� &8  �  �  �"  s    :(� *�� �  8  �  �"    8  �P  �:  ;�4  �  �  <dec �  ;t-  �  <hex �  ;r'  �  ;< �   <oct �  @;� �  �=[)  �   =�%  "�   =�  &�   =dO  )�   =\=  ,�   =�P  /�    =�C  3�   @;zS  6�  �;�O  9�  J=�?  <�  >�  J  ;�7  N  �  ;(  Q  ;�Q  V  ;O  Y   >�9  i�  <in wQ  7  <out zQ   6�� �  �� ?z  �#    /   ?$   �x   �  $,�  -  K  :8   �e  =�  � ?�  "  @�  �4  A("  �J  B."  �A  O�    4"   �A  Q     4"  :"   �A  V0  ;  4"  s    /�
 Y51  �  S  ^  @"  �   /�
 ]�R  �  v  �  @"  �   /� c?  �  �  �  4"  �  �   @_ m.   �  �  4"  �  �   /�3  q89  �  �  �  @"   @.E  ��3  �     4"  �  ."   @�(  ��(  #   .   4"  �   A_Tp 3    �  3ZD  38E  BU  A"  a   �"  s    C9+  N"  �"  s     �� �� �� ?2*  7�   D8   E+  E[  �  [  +  E�  �  8�!   �{  �    ]�  �   \�   �   �D  !�   �3  "�   U>  #�   &�  $�   �  %�   �*  &�    ڡ  '3   $ �U  (3   % TL  )3   & �I  *3   ' Q  +3   ( �C  ,3   ) �J  -3   * 1  .�  , o(  /3   0 �U  03   1 PL  13   2 �I  23   3 Q  33   4 �C  43   5 �J  53   6 F)%  K�  "  s   �   GGT  P"  �   �   s   E3   E�  �  E8   8     E�    s   �  *  �  �  E�  E*  E�  H,   �"  I �  8  E�  E�  �  "  JG   �"  KXF  A�"  K\;  As   LM�T  C"    N\  �"  �"  Oh  �"   d"  Nt  #  #  Oh  �"   J�  2#  LP__p ��    Ja   S#  KXF  N�"  K\;  Ns    N�  a#  v#  Oh  v#  Q__a �{#   p"  L"  e  Nn  �#  �#  Oh  �#   �#  N   �#  �#  Oh  �#  O#  Y"   4"  Nz  �#  �#  Oh  �#  O#  Y"   F"  N  �#  $  Oh  �#  $   :"  N_  $  4$  Oh  �#  Q__a s4$   L"  N�  G$  Q$  Oh  �"   N�  _$  i$  Oh  �"   R�  z$  �$  Oh  �$  O#  Y"   ^"  N  �$  �$  Oh  �$  O#  Y"   j"  S�  ��   ��$  �$  Th  �$  �  �"  N�   �$  %  Oh  %  O#  Y"   �"  U�$  (� ��P   �"%  &  V�$  � W�$  ���! &&  X�$  d_ YQ$  ���! #~%  X_$  d_ Z�"  ��   -X�"  d_   [S#  ���! #Xj#  �_ Xa#  �_ \��    Xj#  �_ Xa#  ` W2#  ���! �&  ]G#  X<#  !` ^�"  ���! V]�"  X�"  !` _�! `�"  6`    a���     b�� U�$  0� ��   �9&  T&  V�$  � a��%  c���+   Nu   b&  w&  Oh  %  K�^  #w&   �"  UT&  R�  �P   ��&  �&  Vb&  � Vk&  �b�b6�aG�,  aP�!,   dU  =�&   �   d�   >�&  dB  ?�&  d�  E�&   �   dB   F�&  dC  G�&  de  H�&  d8  I�&  d�  J�&  d

  XF'   �   d�  YF'  d�
  ZF'  e�   `o'  �   d�  f�'   �   d�  g�'  d�  h�'  d�  n�'   �   d�	  o�'  d�  p�'  dH  v�'   �   d`  w�'  dw  x�'  d   y�'  d~  (   �   d   �(  d�  �(  d  �(  d�   �(  d�  �(  d�	  �(  d�  �`(   �   d  �`(  d  �`(  d�  �`(  d�  ��(   �   d�  ��(  d�  ��(  d�  ��(  dm  ��(     d	  ��(  d2	  ��(  d�  ��(  d9  ��(  d[  �)     dJ  �)  d�  �)  d7  �)  d�  �@)     dI	  �@)  d$	  �@)  d�   �i)   "  dN  �i)  dp  ��)   -  d�  ��)  d:  ��)  d�  )  dd   Æ)  d�  ��)   8  d  ��)  d�  ��)  d�	  ��)   C  d�  ��)  d  �*   N  d�  �*  d�  �*  d�  �*  d+  �B*   Y  d�  �B*  d�   �B*  d  �k*   d  d�
  �k*  d�  �k*  d  �*   o  d   �*  dF  �*  d�  �*   z  d�  ��*  d�  ��*  dD  O�*   �  d�  P�*  d1  Q�*  d�  W+   �  d^  X+  d�  3,+   �  d�  4,+  d�   8I+   �  d�  9I+  dl	  =f+  �  dN  >f+  d^  ?f+  dL  @f+  da  D�+  �  dB  E�+  d�	  F�+  d  G�+  d  H�+  dy  I�+  d�   �+   �  d�  !�+  �  �1  ,  �   f>  Y  !,  �   g  �    �6   ] x� � �V  X"     �� (  _� �7   �  �  8k  �{  k   ]�  k  \�   k  �D  !k  �3  "k  U>  #k  &�  $k  �  %k  �*  &k   ڡ  'q  $�U  (q  %TL  )q  &�I  *q  'Q  +q  (�C  ,q  )�J  -q  *1  .k  ,o(  /q  0�U  0q  1PL  1q  2�I  2q  3Q  3q  4�C  4q  5�J  5q  6 q  �  std # T#  5>   6T#  7�#  @:%  	%  0�=  �n  �b  �q  Fe  �n#  
�3  �=  �  M)  S)   �  eq �<-  Y)    S)  S)   lt ��1  Y)  !  S)  S)   ��  eF  n#  E  `)  `)  n   �K  �9  n  _  `)   �(  
!  `)  �  `)  n  S)   1  �A  f)  �  f)  `)  n   �5  �'  f)  �  f)  `)  n   �3  �A  f)  �  f)  n  �   +  :  �  	  l)   �  �C   �P  �  (  S)   �B  $6  Y)  G  l)  l)   eof (�:  �  ?  ,N0  �  l)    _� �7   �?  �%   K  	\  e%   �e  	_n  �4  	cr)  �J  	dx)  ��  	q�  �  �)   ��  	s�  �  �)  �)   W  	y�  �)  n#    �  �J  
pz  �B  
R  �   %  
k   �B  
A  �)  k  �)    �e  
y�  [V  
k  R  �G  
!   <  
x�  �4  
{�  �J  
|�  �J  
�&  `S  
�)  ~J  
�z  �J  
�  �%  
�  �K  
�R   I  
�R  :!  
��)   %H  
��  �   �3  2k  �G  7{#  t3  B�)  �'  
��O  �)  V  
��N  Y)  [  a  �)   3  
�o+  Y)  x  ~  �)   �P  
��O  �  �  �)   �M  
��P  �  �  �)   �,  
�-  �  �  �)  R   �+  
��R  k  �  �  �)   3  
�   k      �)  �)  �)   �/  !�B  �)  6  R  R  �)   �O  
�|6  I  T  �)  �)    (  ��6  h  s  �)  �)   !�   
�-  k  �  �  �)   "�1  o�*  k  �  �)  �)  R    !�A  
$n%  k  �  �  �)   !�A  
(�I  k  �  �  �)  k   !"A  
,�%  �)      �)   !�1  
2E)  �  -  3  �)   !�/  
6;&  �  K  Q  �)    �>  
:�>  e  k  �)   !S  
A:2  R  �  �  �)  R  u#    �#  
K�(  �  �  �)  R  R  u#   !9  
S>$  R  �  �  �)  R  R   !-U  
[�7  Y)  �    �)  u#   #�5  
d�-  '  k  u#  R   #	1  
m�P  G  k  u#  R   #�3  
v\-  g  k  R  q   #nU  
��-  �  k  �  �   #nU  
�nG  �  k  �  �   #nU  
��   �  k  k  k   #nU  
�IP  �  k  u#  u#   �J  
�rR  n#  	  R  R    �=  ��H  	  /	  �)  R  R  R    V  �)  C	  I	  �)   $�'  
�D*  �)  %�0  
�j	  p	  �)   &�0  ��	  �	  �)  �)   �0  ��	  �	  �)  �)   �0  ��	  �	  �)  �)  R  R   �0  ��	  �	  �)  �)  R  R  �)   �0  �
  
  �)  u#  R  �)   �0  �*
  :
  �)  u#  �)   �0  �J
  _
  �)  R  q  �)   %�0  
"p
  {
  �)  n#   '�  
*,Q  �)  �
  �
  �)  �)   '�  
2�G  �)  �
  �
  �)  u#   '�  
=�%  �)  �
  �
  �)  q   'S� 
f�&  �       �)   'S� 
q�>  �    %  �)   (end 
y<  �  >  D  �)   (end 
�6;  �  ]  c  �)   'I 
��$  �  |  �  �)   'I 
��7  �  �  �  �)   '��  
�lC  �  �  �  �)   '��  
�CM  �  �  �  �)   'r 
��R  R  �  �  �)   '�K  
�r5  R      �)   '�3  
�j=  R  6  <  �)   )�� �  Q  a  �)  R  q   )�� 
��F  v  �  �)  R   'I  
v  R  �  �  �)   )�E  �|U  �  �  �)  R   )�1  
-�  �  �  �)   '�� 
5�?  Y)  �  �  �)   '�:  
D�6  �      �)  R   '�:  
UW  �  7  B  �)  R   (at 
k
/  �  Z  e  �)  R   (at 
��7  �  }  �  �)  R   '�F  
��/  �)  �  �  �)  �)   '�F  
�k:  �)  �  �  �)  u#   '�F  
��H  �)  �  �  �)  q   '@  DA:  �)      �)  �)   '@  U�1  �)  1  F  �)  �)  R  R   '@  )�D  �)  _  o  �)  u#  R   '@  
��*  �)  �  �  �)  u#   '@  �6  �)  �  �  �)  R  q   )�G  
-aN  �  �  �)  q   *�3  �b*  �)  �  �  �)  �)   '�3  
^ 2  �)    -  �)  �)  R  R   '�3  �=  �)  F  V  �)  u#  R   '�3  
z�T  �)  o  z  �)  u#   '�3  
� @  �)  �  �  �)  R  q   )� 
��E  �  �  �)  �  R  q   '� 
�\+  �)  �  �  �)  R  �)   '� 
�u>  �)    )  �)  R  �)  R  R   '� g|=  �)  B  W  �)  R  u#  R   '� 
"�@  �)  p  �  �)  R  u#   '� 
9k<  �)  �  �  �)  R  R  q   '� 
K�'  �  �  �  �)  �  q   'bL  
d�R  �)  �     �)  R  R   'bL  
t�2  �    $  �)  �   'bL  �L&  �  =  M  �)  �  �   '�%  
�9F  �)  f  {  �)  R  R  �)   '�%  
�|<  �)  �  �  �)  R  R  �)  R  R   '�%  ��T  �)  �  �  �)  R  R  u#  R   '�%  
��A  �)  �    �)  R  R  u#   '�%  
b>  �)  -  G  �)  R  R  R  q   '�%  
3%  �)  `  u  �)  �  �  �)   '�%  
'V7  �)  �  �  �)  �  �  u#  R   '�%  
<�+  �)  �  �  �)  �  �  u#   '�%  
Q'S  �)  �  	  �)  �  �  R  q   '�%  
vj.  �)  "  <  �)  �  �  k  k   '�%  
��9  �)  U  o  �)  �  �  u#  u#   '�%  
�C  �)  �  �  �)  �  �  �  �   '�%  
�>/  �)  �  �  �)  �  �  �  �   !�?  ��&  �)  �    �)  R  R  R  q   !�1  �O  �)    9  �)  R  R  u#  R   ,)  
�z-  k  ]  R  q  �)   ++E  �3J  k  �  R  q  �)   '�5  ��)  R  �  �  �)  k  R  R   )n	 @D  �  �  �)  �)   'W�  
�6  u#  �  �  �)   '�A  
%�A  u#      �)   '��  
,Z5  }  %  +  �)   '�(  �;  R  D  Y  �)  u#  R  R   '�(  
I�%  R  r  �  �)  �)  R   '�(  
X�5  R  �  �  �)  u#  R   '�(  �^   R  �  �  �)  q  R   '�(  
v�S  R  �  �  �)  �)  R   '�(  	K  R    +  �)  u#  R  R   '�(  
�o?  R  D  T  �)  u#  R   '�(  J5  R  m  }  �)  q  R   'NW  
��Q  R  �  �  �)  �)  R   'NW  /�I  R  �  �  �)  u#  R  R   'NW  
��,  R  �  �  �)  u#  R   'NW  
��;  R    &  �)  q  R   '�S  
��I  R  ?  O  �)  �)  R   '�S  >T?  R  h  }  �)  u#  R  R   '�S  
05  R  �  �  �)  u#  R   '�S  
$S:  R  �  �  �)  q  R   '�>  
2hL  R  �  �  �)  �)  R   '�>  SUB  R    &  �)  u#  R  R   '�>  
Q�2  R  ?  O  �)  u#  R   '�>  _�K  R  h  x  �)  q  R   '�4  
qT  R  �  �  �)  �)  R   '�4  j�K  R  �  �  �)  u#  R  R   '�4  
��5  R  �  �  �)  u#  R   '�4  N.  R    !  �)  q  R   'U+  
�)  	  :  J  �)  R  R   '��  
�!1  n#  c  n  �)  �)   '��  ��T  n#  �  �  �)  R  R  �)   '��  ��O  n#  �  �  �)  R  R  �)  R  R   '��  �;.  n#  �  �  �)  u#   '��  ��B  n#    &  �)  R  R  u#   '��  ��,  n#  ?  Y  �)  R  R  u#  R     ,!T  q  -�E  �  -�F  �   .�&  .�7  	  �o  >2   �| Cn#  /Q  b�   �  /�F c�  /�R  d�  /3  e�  /�  f�  /�K  g�  /�@  h�   0all i�  ?1�� �d  :!  ��)   NF  �)*  �E  �n  p0  �)*  �%  �5*  2S  �;*  2�R  �;*  23  �;*  2�$  �;*  2�K  �;*  2�@  �;*  2�@  �F*   �4  �Z  �  �  �)    �=  y)  �  �  �)   3�� �    �)  \*  n   3��   %  �)  u#  n   3�� 5  @  �)  n   3N  P  [  �)  n#   3�� k  v  �)  \*    �  �U  �  �  �)  \*   !�&  �.  Y)  �  �  �)    �F  &�;  �  �  �)  b*  �    �9  )�Q  �  �  �)  b*  Q*    WR  ,`2      �)  b*  #*    �S  /=  3  C  �)  #*  /*   4e  7,  S  �)  /*  n    �$  �)   2OD  �)  2gP  �)  2�F  $�)  5< �  6< r�  �.  n    7id �H  �U  �n   2�I  ��)   �  �<?  �  �  *  *   8id �    *  *   9id �&  ,  *   :4H  ��(  n  A  #*    �o  uX  ^  *   �o  ~n  y  *  *   &�o  ��  �  *  u#   �o  ��  �  *  *  u#  �   �o  ��  �  *  *  *  �   5  ��  �  *  n#   *�  ��*  *      *  *   *H�  ��N  7   4  :  *   *U  �9  Y)  R  ]  *  *   *2  �t*  Y)  u  �  *  *   ;jP  �D  �  �  *   <RD  �Q  *  =�o  7�  �  *  �)   >�K  :�N  >�A  =�5  �K  @I  �  �  �    �,  CH<     "   *  *  *  �   �  �     �  � >	  �a  $�   rS  +�#  ?m�  ,e   N   ?��  -e   ?�4  .e   ?;�  /e   ?��  0e   ?� 1e    ?�� 2e   @@b  3e   @�e  4e    @�  5e    ?މ  6e   A�a  �   �.    <s*  =h*  >~*  @+  A+  B3+  CN+  Di+  E�+  F�+  G�+  H�+  ד  ��!  ��  �y  � �k  �4  �r)  ,{�  k   v9,  wi,  {t,  ��,  ��,  ��,  ��,  �-  �--  �B-  �]-  �x-  ��-  ��-  ��-  ��-  ��-  �.  �..  �M.  Rb.  U|.  [�.  \�.  5�+  C#  B��  *��  /  &�F -Q"  k"  =/  C#  /  Y)  n   &�F 9{"  �"  =/  /  Y)  n   C�  E��  q  ("  �"  �"  �0  q   C�  I_�  u#  ("  �"  �"  �0  k  u#   C	�  T}�  q  ("  #  #  �0  q   D	�  X��  u#  ("  2#  �0  k  u#    W�  1C/  ("   E)%  Kk  n#  n#  u#   Fint {#  q  GGT  P�#  >   �  �#  �  �  o  �	  �  qW  !n#    "�#  �  #  .  <�#  `  Dn#  �  W�#  �  _�#  �  en#  t   mn#  a  un#    ~n#  �  �n#  3  �n#  �  �n#  H  �n#  y  �n#    �n#  s  �n#  T   �n#  �  �n#  F  �n#  �  �n#  �  �n#    �n#  V  �n#  �  Hs  N�#  �  V�#  \	  2n#  o  7n#  �  <n#  �  Cn#  �  n#  1%  IJpO qO !2%  K$   E%)  	�  $,n  -y  K  :�&  �e  =n  � ?k  "  @u#  �4  Ar)  �J  Bx)  �A  O�%  �%  ~)   �A  Q�%  �%  ~)  �)   �A  V�%  �%  ~)  n#   *�
 Y51  }%  &  &  �)  �%   *�
 ]�R  �%  4&  ?&  �)  �%   *� c?  }%  W&  g&  ~)  q%  +%   L_ m.   {&  �&  ~)  }%  q%   *�3  q89  q%  �&  �&  �)   L.E  ��3  �&  �&  ~)  }%  x)   L�(  ��(  �&  �&  ~)  }%   M_Tp q   e%  NZD  �)  OF�  �k   P��  �U!  P�4  �k!  P� �`!  %��  �N'  T'  �+   Q��  �e'  p'  �+  �+   '*  ��}  #'  �'  �'  ,   'Ư  �?s  0'  �'  �'  ,   '�F  �Ϭ  ,  �'  �'  �+   '�F  ��  �&  �'  �'  �+  n#   'a�  �
�  ,  
(  (  �+   'a�   ��  �&  )(  4(  �+  n#   '�:  ,�  #'  M(  X(  ,  '   '�F  		n  ,  q(  |(  �+  '   '(*  ��  �&  �(  �(  ,  '   ' I  h�  ,  �(  �(  �+  '   '�O  7k  �&  �(  �(  ,  '   'WC  ]�  �+  )  )  ,   ,{�  k  ,�  	   .8E  �&   �� �� �� K2*  7M)  R8�   S�  S�  �  �  �  S	  Sq  S{#  e%  S�&  �&  �  S  �)    �   n#    �  	    S  S�  S	  T7   �)  U Y    �)   *  u#  �  S2   2   �  S"   "   /*  '   k  T#*  F*  U TQ*  Q*  U W*  #*  S,   ,   �l  %   j�  #%   Vtm ,,+  ,g  .n#   �  /n#  �  0n#  ��  1n#  ��  2n#  ��  3n#  ��  4n#  �  5n#  d�  6n#   ��  7%   $~�  8u#  ( G\�  >s*  Eѯ  H,)  3+  h*  h*   E��  Mh*  H+  H+   ~*  E�  Ch*  c+  c+   h*  E#�  ak  ~+  ~+   �+  ~*  E�� fk  �+  �+   �+  h*  E��  WH+  �+  �+   E[v  \H+  �+  �+   E��  R,   �+  k  ,   u#  ~+   �&  S,  k  )  S�&  W *  9,  �   n#   Xrem  n#   +    ,  W #@  i,  �   $%    Xrem  %%    A   &D,  E�  �n#  �,  �,   �,  YE�   >,)  �,  u#   E�   Hn#  �,  u#   E�   I%   �,  u#   E�   ��$  �,  +%  +%  ,   ,   �,   �,  Zn#  -  +%  +%   [div  9,  --  n#  n#   E     �k  B-  u#   \�    i,  ]-  %   %    \�   .n#  x-  u#  ,    \�   \,   �-  �)  u#  ,    \3   >n#  �-  �)  u#  ,    ]�   �-  �$  ,   ,   �,   Gk�  qn#  ^�   |�-  �#   E   W,)  .  u#  5*   E   f%   ..  u#  5*  n#   E�   g7   M.  u#  5*  n#   E?   �n#  b.  u#   E��  !En#  |.  u#  u#   E��  !Uk  �.  n#   E��  !Ok  �.  k  u#   E��  !F,   �.  k  u#  ,    �  _�  �.  �.  `h  �.  a4&  rn   �.  B   b�   $/  /  `h  /   �.  e   c1"  d$/  ��  P�   �("  n#  _A"   W/  �/  `h  �/  C#  ep� -/  e(� -Y)  e4&  .n   =/  fI/  E� `��   ��/  �/  gW/  V` h`/  �ge/  u` gp/  �` g{/  �` i�.  a�" 1g�.  �` g�.  �`   _k"   0  /0  `h  �/  ep� 9/  e(� 9Y)  e4&  9n   f�/  .�  ��   �J0  �0  g0  �` g0  a g0  /a g#0  Ca i�.  �8" <g�.  Wa g�.  ka   N#  j�"  ��   ��0  �0  kh  �0  � l__c Eq  �m���6   �0  j�"  ��A   ��0  !1  kh  �0  � n�a  Ik  �a o�a  Iu#  �m���6   j�"  �   �81  \1  kh  �0  � l__c Tq  �m��6   j#  0�A   �s1  �1  kh  �0  � n�a  Xk  �a o�a  Xu#  �m_��6   pU  =�1   �#  p�   >�1  pB  ?�1  p�  E�1   �#  pB   F�1  pC  G�1  pe  H�1  p8  I�1  p�  J�1  p

  X(2   �#  p�  Y(2  p�
  Z(2  q�   `Q2  $  p�  fb2   $  p�  gb2  p�  hb2  p�  n�2   $  p�	  o�2  p�  p�2  pH  v�2   %$  p`  w�2  pw  x�2  p   y�2  p~  �2   0$  p   ��2  p�  ��2  p  ��2  p�   ��2  p�  ��2  p�	  ��2  p�  �B3   ;$  p  �B3  p  �B3  p�  �B3  p�  �w3   F$  p�  �w3  p�  �w3  p�  �w3  pm  ��3   Q$  p	  ��3  p2	  ��3  p�  ��3  p9  ��3  p[  ��3   \$  pJ  ��3  p�  ��3  p7  ��3  p�  �"4   g$  pI	  �"4  p$	  �"4  p�   �K4   r$  pN  �K4  pp  �h4   }$  p�  �h4  p:  �h4  p�  �h4  pd   �h4  p�  ɩ4   �$  p  ʩ4  p�  ˩4  p�	  ��4   �$  p�  ��4  p  ��4   �$  p�  ��4  p�  ��4  p�  ��4  p+  �$5   �$  p�  �$5  p�   �$5  p  �M5   �$  p�
  �M5  p�  �M5  p  �v5   �$  p   �v5  pF  �v5  p�  �5   �$  p�  ��5  p�  ��5  pD  O�5   �$  p�  P�5  p1  Q�5  p�  W�5   �$  p^  X�5  p�  36   �$  p�  46  p�   8+6   �$  p�  9+6  pl	  =H6  
%  pN  >H6  p^  ?H6  pL  @H6  pa  D}6  %  pB  E}6  p�	  F}6  p  G}6  p  H}6  py  I}6  p�   �6    %  p�  !�6  Ek�  "�n#  �6  n#   r��  "�n#  n#    �   � w� ^� �V  �"     �� (  _� �7   �  �  8k  �{  k   ]�  k  \�   k  �D  !k  �3  "k  U>  #k  &�  $k  �  %k  �*  &k   ڡ  'q  $�U  (q  %TL  )q  &�I  *q  'Q  +q  (�C  ,q  )�J  -q  *1  .k  ,o(  /q  0�U  0q  1PL  1q  2�I  2q  3Q  3q  4�C  4q  5�J  5q  6 q  �  std  �  5>   6�  7�  @w  	%  0_� �7   �?  �%   <�  =�  >�  @  A�  B�  C�  D�  E�  F  G/  HD  Rh  U�  [�  \�  
_}  �  ��  *��  �  M  ]  �  �  �    ~  3��  �  u  �  �  k  �  �   !T  q   ,   )%  Kk  �  �  �   int �  q  GT  P�  >   �  	�  �  �  o  �	  �  qW  	!�    	"  �  #  .  
<  `  
D�  �  
W  �  
_  �  
e�  t   
m�  a  
u�    
~�  �  
��  3  
��  �  
��  H  
��  y  
��    
��  s  
��  T   
ȴ  �  
д  F  
״  �  
�  �  
�    
�  V  
�  �  s  N�  �  V�  \	  2�  o  7�  �  <�  �  C�  �  �  pO qO !o  $   E�  	�  $,�  -�   �� �� �� 2*  7�  8�   �    �l  %   j�  #%   tm ,,  ,g  .�   �  /�  �  0�  ��  1�  ��  2�  ��  3�  ��  4�  �  5�  d�  6�   ��  7%   $~�  8�  ( \�  >�  ѯ  H�  �  �  �   ��  M�  �  �   �  �  C�  �  �   �  #�  ak  �  �   �  �  �� fk         �  ��  W�  /     [v  \�  D     ��  R,   h  k  ,   �  �   ��  E�  �  �  �   ��  Uk  �  �   ��  Ok  �  k  �   ��  F,   �  k  �  ,    �  5  ��    ��  4  h  4  � ��  *�  ���  +�  ��" q� -�  �a ��h    �  ]  ��   �P  �  h  4  b "y  3k  b DK 3�  >b __n 4�  � ���  !��  "U  
=�   )  "�   
>�  "B  
?�  "�  
E�   4  "B   
F�  "C  
G�  "e  
H�  "8  
I�  "�  
J�  "

  
X   ?  "�  
Y  "�
  
Z  #�   
`G  J  "�  
fX   U  "�  
gX  "�  
hX  "�  
n�   `  "�	  
o�  "�  
p�  "H  
v�   k  "`  
w�  "w  
x�  "   
y�  "~  
�   v  "   
��  "�  
��  "  
��  "�   
��  "�  
��  "�	  
��  "�  
�8	   �  "  
�8	  "  
�8	  "�  
�8	  "�  
�m	   �  "�  
�m	  "�  
�m	  "�  
�m	  "m  
��	   �  "	  
��	  "2	  
��	  "�  
��	  "9  
��	  "[  
��	   �  "J  
��	  "�  
��	  "7  
��	  "�  
�
   �  "I	  
�
  "$	  
�
  "�   
�A
   �  "N  
�A
  "p  
�^
   �  "�  
�^
  ":  
�^
  "�  
�^
  "d   
�^
  "�  
ɟ
   �  "  
ʟ
  "�  
˟
  "�	  
��
   �  "�  
��
  "  
��
   �  "�  
��
  "�  
��
  "�  
��
  "+  
�   �  "�  
�  "�   
�  "  
�C   �  "�
  
�C  "�  
�C  "  
�l     "   
�l  "F  
�l  "�  
�     "�  
��  "�  
��  "D  O�   "  "�  P�  "1  Q�  "�  W�   -  "^  X�  "�  3   8  "�  4  "�   8!   C  "�  9!  "l	  =>  N  "N  >>  "^  ?>  "L  @>  "a  Ds  Y  "B  Es  "�	  Fs  "  Gs  "  Hs  "y  Is  "�   �   d  "�  !�      h H� 
� �V  ϰ (  _� �/   �  �  �  H   �  �  o  �	  pW   o   �  qW  !�   int   "�   �    #�   #  Fd v   .  <v   `  D�   �  Wv   �  _�   �  e�   t   m�   a  u�     ~�   �  ��   3  ��   �  ��   H  ��   y  ��     ��   s  ��   T   ȁ   �  Ё   F  ׁ   �  ��   �  �     �   V  �   6   �  s  N=   �  V=   \	  2�   o  7�   �  <�   �  C�   �  �   =   	\  �   gX  �   X\  &+  X\  X,@  	$Z  .�    	\ /=   	� 1  	Z  2$   	K]  3=   	�_  4$   	\W  5$   	�Z  6$   	-_  8_   	VY  9�  $	`  :�  (	�Y  ;�  ,	7_  <�  0	BY  =�  4	b\  >�  8	\  ?�  <	7Y  @�  @	 Z  A	  D	SX  B	  H	n4 Dd   L	`  FY  P	*5 GY  T 
  Y  �  $   Y   +  @  
  ~  ~  $   Y   �  e  
�   �  Y  
  �    �  

  �  Y   �  
�   �  Y   �  
Y  �  �  �  Y   �  6   �  	  Y   �  	pO qO 	!  std  }  @  %  0_� 
�/   5�  6�  7  �?  
�   b   c,  e7  fO  gd  hz  i�  j�  k�  l�  m�  q  r;  tZ  uz  v�  x�  y�  |�  ~�  ��  �	  �.	  �@	  �V	  �z	  ��	  ��	  �� 4�  cin 8T�  *  ִ 6�  ��  9��  D  M�  :H�  D  A�  ;<�  D   $   ��  �  $,;  -[   �� �� �� 2*  7�  84   �  �  8�  	�{  �   	]�  �  	\�   �  	�D  !�  	�3  "�  	U>  #�  	&�  $�  	�  %�  	�*  &�   	ڡ  '6   $	�U  (6   %	TL  )6   &	�I  *6   '	Q  +6   (	�C  ,6   )	�J  -6   *	1  .�  ,	o(  /6   0	�U  06   1	PL  16   2	�I  26   3	Q  36   4	�C  46   5	�J  56   6 )%  K�    �   �   GT  P  �    �^  !
  Z  1I  I      aY  ��   d  I   \  C�   z  I   xZ  M�   �  I   `  ��   �  I   �^  r�   �  I   _X  ��   �  I  �   ,  �_  ��  �  �  �   I   �\  �I    �  �   4Z  �$   ;  ~  $   $   I   7`  �I  Z  �  �  I   >]  	�   z  I     �    �Z  �   �  I  �   �  ,  �Y      �  I   �Y  ��   �  I   \  ��   �_  0�  �  �   �]  W�  �   D[  T�   	  �   �[  a�   .	  �  �   �\  )@	  I   Y@ �V	  I  �   �[     z	  I  �  �   $    �]  iI  D]  w�  �	  �   }W  ��   �	  �   I   ��  L?
  M"  N}  � Rt  %�  T�  �	  ��  U@�  �	  ��  V�  �	  � X�  ?�  Z��  
  ��  [3�  
  ��  \��  
   U  =K
   �   �   >K
  B  ?K
  �  Et
   �   B   Ft
  C  Gt
  e  Ht
  8  It
  �  Jt
  

  X�
   �   �  Y�
  �
  Z�
  �   `�
  �   �  f�
   �   �  g�
  �  h�
  �  n$   �   �	  o$  �  p$  H  vM   �   `  wM  w  xM     yM  ~  �        ��  �  ��    ��  �   ��  �  ��  �	  ��  �  ��       ��    ��  �  ��  �  �     �  �  �  �  �  �  m  �E   $  	  �E  2	  �E  �  �E  9  �E  [  ��   /  J  ��  �  ��  7  ��  �  ��   :  I	  ��  $	  ��  �   ��   E  N  ��  p  �   P  �  �  :  �  �  �  d   �  �  �B   [    �B  �  �B  �	  �k   f  �  �k    ؈   q  �  و  �  ڈ  �  ۈ  +  �   |  �  �  �   �    ��   �  �
  ��  �  ��    �   �     �  F  �  �  �8   �  �  �8  �  �8  D  Oa   �  �  Pa  1  Qa  �  W�   �  ^  X�  �  3�   �  �  4�  �   8�   �  �  9�  l	  =�  �  N  >�  ^  ?�  L  @�  a  D  �  B  E  �	  F    G    H  y  I  �   c   �  �  !c  6   �   �  ' !�	  �W!�	  �W!�	  `W6   �   �  _ !
   W! 
  �V!/
   V6   �   �  � !5  �Z6      �  � !O  �Y!^   Y!m  @X �   
 � ҵ �V  (#     r� (  �  �  �  E   �  �  o  �	  �  qW  !s   int   "�   �  #  .  <h   `  Ds   �  Wh   �  _z   �  es   t   ms   a  us     ~s   �  �s   3  �s   �  �s   H  �s   y  �s     �s   s  �s   T   �s   �  �s   F  �s   �  �s   �  �s     �s   V  �s   3   �  s  N:   �  V:   \	  2s   o  7s   �  <s   �  Cs   �  	s   �  �  3   	
pO qO 
!�  
std  �  @�  5�  6�  7�  %  0�=  ��  �b  �3   Fe  �s   �3  �=  p  E  K   @  eq �<-  Q  �  K  K   lt ��1  Q  �  K  K   ��  eF  s   �  X  X  �   �K  �9  �  �  X   �(  
!  X    X  �  K   1  �A  ^  5  ^  X  �   �5  �'  ^  Y  ^  X  �   �3  �A  ^  }  ^  �  @   +  :  @  �  d   K  �C   �P  K  �  K   �B  $6  Q  �  d  d   eof (�:  K  ?  ,N0  K  d    _� �,   �?  �%   �8  �  �@  ]  0  @  �  s   |   �  TP  e  �  s   |  \	   {'  E8  �  ��  �  �  s   |   !T  3   �E  4   �Y  8  �% g�  �  �  �  s   |   ̾ ]�  �  �  s   |  �
   {'  E8  ̾ ^  %  �  s   |   !T  3   �E  4   �M  T  !T  3   �E  4   `'  �w  �>  �3    !T  3    $ ��    �      l* 4�  �  v  s   |  �   !k* ;w  �  �  v  s   |   l* >�    v  s   |   !T  3   �E  4   �E  �  !`V    5  @  �  s    aV  �Q  W  �   !T  3   �E  4  "i3 ~P4  y  �  �    #�� ��� T  !T  3   3     �  8�  $�{  �   $]�  �  $\�   �  $�D  !�  $�3  "�  $U>  #�  $&�  $�  $�  %�  $�*  &�   $ڡ  '3   $$�U  (3   %$TL  )3   &$�I  *3   '$Q  +3   ($�C  ,3   )$�J  -3   *$1  .�  ,$o(  /3   0$�U  03   1$PL  13   2$�I  23   3$Q  33   4$�C  43   5$�J  53   6 %)%  K�  �  s   �   &GT  P�  �  '$   '  �  $,�  -   �� �� �� '2*  7E  (8-   )@  )p  �  p  @  )�    s   w  �  8    *  �  �  +h  �  +#  q   �    *  �  �  +h  �  +#  q  +�!  �   �  |  �  *�  	  	  +h  	  +#  q  +�!  #	   �  |  *�  6	  R	  +h  R	  +#  q  +�!  W	   v  |  e  *@  p	  �	  +h  �  +#  q  +�!  �	  ,(  T\	   |  *@  �	  �	  +h  �   *q  �	  �	  +h  �  +#  q  +�!  �	   |  -(	  �� ��   ��	  '
  .6	  ]b /�  ��   ;.�  ~b 0��  -(	  �  �%   �B
  �
  16	  � 2(	  �   ;�
  .6	  �b /�  �   ;.�  �b 3�  4%��   5�  P�   ��
  !T  3   6__c �3   � �  *�  �
  �
  +h  	  +#  q  +�!  �
  ,(  ]�
   |  *�  
  2  +h  R	  +#  q  +�!  2  7(  4�   |  -�
  � `��   �R    1
  � 1  �1%  �2�
  r�!   5�  .�
  �b .�
  3c .�
  uc 8��i   9b	  ���" 5�  .�	  �c .�	  �c .p	  #d 8��i   2�  ��   5  1	  v�1	  S 8���   -�
  Y� ���   �&  �  1
  � 1%  �2�	  ��F   5Y  .�	  ed 3� 2�
  E�   5�  .�
  �d 1�
  L	�.�
  �d 8b�i   9b	  d��" 5�  .�	  (e :�	  .p	  Se 8y�i   2�  ��   5�  1�  s�3�� 8���   -(	  � ��<   �  u  16	  � 1H	  �2�  ��   ;O  1�  �#�1�  � #� /�  ��   ;1	  �#�1	  �   *  �  �  +h  	  +#  q  +�!  �   |  *�  �  �  +h  R	  +#  q  +�!  �   |  -�  ��  ��   ��  �  1�  � 1�  �2u  �%   ?.  .�  �e .�  �e 80�i   9�	  0��" ?^  .�	   f .�	  Bf 8L�i   2�  i�   ?�  1	  v�1	  S 8���   -�  O� ���   ��  _  1�  � 2�	  ��F   ?�  .�	  �f 3�� 2u  ��    ?  1�  L	�.�  �f 8��i   9�	  ��# ?2  :�	  .�	  g 8�i   2�  )�   ?U  1�  s�39� 8A��   ;U  =k   �   ;�   >k  ;B  ?k  ;�  E�   �   ;B   F�  ;C  G�  ;e  H�  ;8  I�  ;�  J�  ;

  X�   �   ;�  Y�  ;�
  Z�  <�   `
  �   ;�  f   �   ;�  g  ;�  h  ;�  nD   �   ;�	  oD  ;�  pD  ;H  vm   �   ;`  wm  ;w  xm  ;   ym  ;~  �   �   ;   ��  ;�  ��  ;  ��  ;�   ��  ;�  ��  ;�	  ��  ;�  ��   �   ;  ��  ;  ��  ;�  ��  ;�  �0   �   ;�  �0  ;�  �0  ;�  �0  ;m  �e     ;	  �e  ;2	  �e  ;�  �e  ;9  �e  ;[  ��     ;J  ��  ;�  ��  ;7  ��  ;�  ��     ;I	  ��  ;$	  ��  ;�   �   "  ;N  �  ;p  �!   -  ;�  �!  ;:  �!  ;�  �!  ;d   �!  ;�  �b   8  ;  �b  ;�  �b  ;�	  ы   C  ;�  ҋ  ;  ب   N  ;�  ٨  ;�  ڨ  ;�  ۨ  ;+  ��   Y  ;�  ��  ;�   ��  ;  �   d  ;�
  �  ;�  �  ;  �/   o  ;   �/  ;F  �/  ;�  �X   z  ;�  �X  ;�  �X  ;D  O�   �  ;�  P�  ;1  Q�  ;�  W�   �  ;^  X�  ;�  3�   �  ;�  4�  ;�   8�   �  ;�  9�  ;l	  =  �  ;N  >  ;^  ?  ;L  @  ;a  D6  �  ;B  E6  ;�	  F6  ;  G6  ;  H6  ;y  I6  ;�  	 �   �  ;�  	!�  �  �1  �  �   =>  Y  �    21   x ̶ �� �V  �#     #� (  _� �7   �  �  8k  �{  k   ]�  k  \�   k  �D  !k  �3  "k  U>  #k  &�  $k  �  %k  �*  &k   ڡ  'q  $�U  (q  %TL  )q  &�I  *q  'Q  +q  (�C  ,q  )�J  -q  *1  .k  ,o(  /q  0�U  0q  1PL  1q  2�I  2q  3Q  3q  4�C  4q  5�J  5q  6 q  �  std  Y!  5>   6Y!  7�!  @?#  	%  0�=  �n  �b  �q  Fe  �s!  
�3  �=  �  R'  X'   �  eq �<-  ^'    X'  X'   lt ��1  ^'  !  X'  X'   ��  eF  s!  E  e'  e'  n   �K  �9  n  _  e'   �(  
!  e'  �  e'  n  X'   1  �A  k'  �  k'  e'  n   �5  �'  k'  �  k'  e'  n   �3  �A  k'  �  k'  n  �   +  :  �  	  q'   �  �C   �P  �  (  X'   �B  $6  ^'  G  q'  q'   eof (�:  �  ?  ,N0  �  q'    _� 	�7   �?  	�%   K  
\  j#   �e  
_n  �4  
cw'  �J  
d}'  ��  
q�  �  �'   ��  
s�  �  �'  �'   W  
y�  �'  s!    �  �J  pz  �B  R  �   %  k   �B  A  �'  k  �'    �e  y�  [V  k  R  �G  !   <  x�  �4  {�  �J  |�  �J   %  `S  �'  ~J  �z  �J  �  �%  �  �K  �R   I  �R  :!  ��'   %H  ��  �   �3  2k  �G  7�!  t3  B�'  �'  ��O  �'  V  ��N  ^'  [  a  �'   3  �o+  ^'  x  ~  �'   �P  ��O  �  �  �'   �M  ��P  �  �  �'   �,  �-  �  �  �'  R   �+  ��R  k  �  �  �'   3  �   k      �'  �'  �'   �/  !�B  �'  6  R  R  �'   �O  �|6  I  T  �'  �'    (  ��6  h  s  �'  �'   !�   �-  k  �  �  �'   "�1  o�*  k  �  �'  �'  R    !�A  $n%  k  �  �  �'   !�A  (�I  k  �  �  �'  k   !"A  ,�%  �'      �'   !�1  2E)  �  -  3  �'   !�/  6;&  �  K  Q  �'    �>  :�>  e  k  �'   !S  A:2  R  �  �  �'  R  z!    �#  K�(  �  �  �'  R  R  z!   !9  S>$  R  �  �  �'  R  R   !-U  [�7  ^'  �    �'  z!   #�5  d�-  '  k  z!  R   #	1  m�P  G  k  z!  R   #�3  v\-  g  k  R  q   #nU  ��-  �  k  �  �   #nU  �nG  �  k  �  �   #nU  ��   �  k  k  k   #nU  �IP  �  k  z!  z!   �J  �rR  s!  	  R  R    �=  ��H  	  /	  �'  R  R  R    V  �)  C	  I	  �'   $�'  �D*  �'  %�0  �j	  p	  �'   &�0  ��	  �	  �'  �'   �0  ��	  �	  �'  �'   �0  ��	  �	  �'  �'  R  R   �0  ��	  �	  �'  �'  R  R  �'   �0  �
  
  �'  z!  R  �'   �0  �*
  :
  �'  z!  �'   �0  �J
  _
  �'  R  q  �'   %�0  "p
  {
  �'  s!   '�  *,Q  �'  �
  �
  �'  �'   '�  2�G  �'  �
  �
  �'  z!   '�  =�%  �'  �
  �
  �'  q   'S� f�&  �       �'   'S� q�>  �    %  �'   (end y<  �  >  D  �'   (end �6;  �  ]  c  �'   'I ��$  �  |  �  �'   'I ��7  �  �  �  �'   '��  �lC  �  �  �  �'   '��  �CM  �  �  �  �'   'r ��R  R  �  �  �'   '�K  �r5  R      �'   '�3  �j=  R  6  <  �'   )�� �  Q  a  �'  R  q   )�� ��F  v  �  �'  R   'I  v  R  �  �  �'   )�E  �|U  �  �  �'  R   )�1  -�  �  �  �'   '�� 5�?  ^'  �  �  �'   '�:  D�6  �      �'  R   '�:  UW  �  7  B  �'  R   (at k
/  �  Z  e  �'  R   (at ��7  �  }  �  �'  R   '�F  ��/  �'  �  �  �'  �'   '�F  �k:  �'  �  �  �'  z!   '�F  ��H  �'  �  �  �'  q   '@  DA:  �'      �'  �'   '@  U�1  �'  1  F  �'  �'  R  R   '@  )�D  �'  _  o  �'  z!  R   '@  ��*  �'  �  �  �'  z!   '@  �6  �'  �  �  �'  R  q   )�G  -aN  �  �  �'  q   *�3  �b*  �'  �  �  �'  �'   '�3  ^ 2  �'    -  �'  �'  R  R   '�3  �=  �'  F  V  �'  z!  R   '�3  z�T  �'  o  z  �'  z!   '�3  � @  �'  �  �  �'  R  q   )� ��E  �  �  �'  �  R  q   '� �\+  �'  �  �  �'  R  �'   '� �u>  �'    )  �'  R  �'  R  R   '� g|=  �'  B  W  �'  R  z!  R   '� "�@  �'  p  �  �'  R  z!   '� 9k<  �'  �  �  �'  R  R  q   '� K�'  �  �  �  �'  �  q   'bL  d�R  �'  �     �'  R  R   'bL  t�2  �    $  �'  �   'bL  �L&  �  =  M  �'  �  �   '�%  �9F  �'  f  {  �'  R  R  �'   '�%  �|<  �'  �  �  �'  R  R  �'  R  R   '�%  ��T  �'  �  �  �'  R  R  z!  R   '�%  ��A  �'  �    �'  R  R  z!   '�%  b>  �'  -  G  �'  R  R  R  q   '�%  3%  �'  `  u  �'  �  �  �'   '�%  'V7  �'  �  �  �'  �  �  z!  R   '�%  <�+  �'  �  �  �'  �  �  z!   '�%  Q'S  �'  �  	  �'  �  �  R  q   '�%  vj.  �'  "  <  �'  �  �  k  k   '�%  ��9  �'  U  o  �'  �  �  z!  z!   '�%  �C  �'  �  �  �'  �  �  �  �   '�%  �>/  �'  �  �  �'  �  �  �  �   !�?  ��&  �'  �    �'  R  R  R  q   !�1  �O  �'    9  �'  R  R  z!  R   ,)  �z-  k  ]  R  q  �'   ++E  �3J  k  �  R  q  �'   '�5  ��)  R  �  �  �'  k  R  R   )n	 @D  �  �  �'  �'   'W�  �6  z!  �  �  �'   '�A  %�A  z!      �'   '��  ,Z5  }  %  +  �'   '�(  �;  R  D  Y  �'  z!  R  R   '�(  I�%  R  r  �  �'  �'  R   '�(  X�5  R  �  �  �'  z!  R   '�(  �^   R  �  �  �'  q  R   '�(  v�S  R  �  �  �'  �'  R   '�(  	K  R    +  �'  z!  R  R   '�(  �o?  R  D  T  �'  z!  R   '�(  J5  R  m  }  �'  q  R   'NW  ��Q  R  �  �  �'  �'  R   'NW  /�I  R  �  �  �'  z!  R  R   'NW  ��,  R  �  �  �'  z!  R   'NW  ��;  R    &  �'  q  R   '�S  ��I  R  ?  O  �'  �'  R   '�S  >T?  R  h  }  �'  z!  R  R   '�S  05  R  �  �  �'  z!  R   '�S  $S:  R  �  �  �'  q  R   '�>  2hL  R  �  �  �'  �'  R   '�>  SUB  R    &  �'  z!  R  R   '�>  Q�2  R  ?  O  �'  z!  R   '�>  _�K  R  h  x  �'  q  R   '�4  qT  R  �  �  �'  �'  R   '�4  j�K  R  �  �  �'  z!  R  R   '�4  ��5  R  �  �  �'  z!  R   '�4  N.  R    !  �'  q  R   'U+  �)  	  :  J  �'  R  R   '��  �!1  s!  c  n  �'  �'   '��  ��T  s!  �  �  �'  R  R  �'   '��  ��O  s!  �  �  �'  R  R  �'  R  R   '��  �;.  s!  �  �  �'  z!   '��  ��B  s!    &  �'  R  R  z!   '��  ��,  s!  ?  Y  �'  R  R  z!  R     ,!T  q  -�E  �  -�F  �   .�&  .�7  	  �o  >2   �| Cs!  /Q  b�   �  /�F c�  /�R  d�  /3  e�  /�  f�  /�K  g�  /�@  h�   0all i�  ?1�� �d  :!  ��'   NF  �-(  �E  �n  p0  �-(  �%  �9(  2S  �?(  2�R  �?(  23  �?(  2�$  �?(  2�K  �?(  2�@  �?(  2�@  �J(   �4  �Z  �  �  �'    �=  y)  �  �  �'   3�� �    �'  `(  n   3��   %  �'  z!  n   3�� 5  @  �'  n   3N  P  [  �'  s!   3�� k  v  �'  `(    �  �U  �  �  �'  `(   !�&  �.  ^'  �  �  �'    �F  &�;  �  �  �'  f(  �    �9  )�Q  �  �  �'  f(  U(    WR  ,`2      �'  f(  '(    �S  /=  3  C  �'  '(  3(   4e  7,  S  �'  3(  n    �$  �'   2OD  �'  2gP  �'  2�F  $�'  5< �  6< r�  *  n    7id �H  �U  �n   2�I  ��'   �  �<?  �  �  (  !(   8id �    (  !(   9id �&  ,  (   :4H  ��(  n  A  '(    �o  uX  ^  	(   �o  ~n  y  	(  (   &�o  ��  �  	(  z!   �o  ��  �  	(  (  z!  �   �o  ��  �  	(  (  (  �   5  ��  �  	(  s!   *�  ��*  (      	(  (   *H�  ��N  7   4  :  (   *U  �9  ^'  R  ]  (  (   *2  �t*  ^'  u  �  (  (   ;jP  �D  �  �  (   <RD  �Q  (  =�o  7�  �  	(  �'   >�K  :�N  >�A  =�5  �K  @I  �  �  �    �,  CH<     "   	(  (  (  �   �  �     �  � >	  <w(  =l(  >�(  @)  A)  B7)  CR)  Dm)  E�)  F�)  G�)  H�)  ד  ��   ��  �y  � �k  �4  �w'  ,{�  k   ?0T  �   3��  :�   �   G*  n   ,!T  q   5�N  M!  @��  '��  !  #!  v*  M!   A�o  A�   8!  C!  v*  s!   ,!T  q   W�  1|*   B)%  Kk  s!  s!  z!   Cint �!  q  DGT  P�!  >   �  �!  �  �  o  �	  �  qW  !s!    "�!  �  #  .  <�!  `  Ds!  �  W�!  �  _�!  �  es!  t   ms!  a  us!    ~s!  �  �s!  3  �s!  �  �s!  H  �s!  y  �s!    �s!  s  �s!  T   �s!  �  �s!  F  �s!  �  �s!  �  �s!    �s!  V  �s!  �  Es  N�!  �  V�!  \	  2s!  o  7s!  �  <s!  �  Cs!  �  s!  6#  FGpO qO !7#  H$   E*'  	�  $,n  -y  K  :�$  �e  =n  � ?k  "  @z!  �4  Aw'  �J  B}'  �A  O�#  �#  �'   �A  Q�#  �#  �'  �'   �A  V�#  �#  �'  s!   *�
 Y51  �#  $  !$  �'  �#   *�
 ]�R  �#  9$  D$  �'  �#   *� c?  �#  \$  l$  �'  v#  0#   @_ m.   �$  �$  �'  �#  v#   *�3  q89  v#  �$  �$  �'   @.E  ��3  �$  �$  �'  �#  }'   @�(  ��(  �$  �$  �'  �#   I_Tp q   j#  JZD  �'  KF�  �k   L��  ��   L�4  ��   L� ��   %��  �S%  Y%  �)   M��  �j%  u%  �)  *   '*  ��}  (%  �%  �%  *   'Ư  �?s  5%  �%  �%  *   '�F  �Ϭ  *  �%  �%  �)   '�F  ��   %  �%  �%  �)  s!   'a�  �
�  *  &  &  �)   'a�   ��   %  .&  9&  �)  s!   '�:  ,�  (%  R&  ]&  *  %   '�F  		n  *  v&  �&  �)  %   '(*  ��   %  �&  �&  *  %   ' I  h�  *  �&  �&  �)  %   '�O  7k   %  �&  �&  *  %   'WC  ]�  *  '  '  *   ,{�  k  ,�  	   .8E   %   �� �� �� H2*  7R'  N8�   O�  O�  �  �  �  O	  Oq  O�!  j#  O�$  �$  �  O    �   s!  s!    �  	    O  O�  O	  P7   �'  Q Y    �'  (  z!  �  O2   2   �  O"   "   3(  '   k  P'(  J(  Q PU(  U(  Q [(  '(  O,   ,   �l  %   j�  #%   Rtm ,,)  ,g  .s!   �  /s!  �  0s!  ��  1s!  ��  2s!  ��  3s!  ��  4s!  �  5s!  d�  6s!   ��  7%   $~�  8z!  ( D\�  >w(  Bѯ  H1'  7)  l(  l(   B��  Ml(  L)  L)   �(  B�  Cl(  g)  g)   l(  B#�  ak  �)  �)   �)  �(  B�� fk  �)  �)   �)  l(  B��  WL)  �)  �)   B[v  \L)  �)  �)   B��  R,   �)  k  ,   z!  �)    %  O*  k  $'  O %  �  S�  ,*  B*  Th  B*  U4&  rn   *  �   S�   [*  q*  Th  q*  U4&  :n   G*  �   s!  V!  P��   ��*  0+  Wh  0+  � XM!  �Y��)   �*  Z__i 4n  :g  Y��   �*  Z__i 7n  Yg  [M*  ��G   +&+  \d*   ][*  P^*  ��   ?\5*   ],*  P  _���0   v*  S#!   C+  V+  Th  0+  T#  �'   `5+  _� P�B   �q+  �+  ]C+  � a�b��_��1   c5+  �� ��   ��+  �+  ]C+  � _��V+  d��$1   eU  =�+   �!  e�   >�+  eB  ?�+  e�  E�+   �!  eB   F�+  eC  G�+  ee  H�+  e8  I�+  e�  J�+  e

  XE,   �!  e�  YE,  e�
  ZE,  f�   `n,  	"  e�  f,   "  e�  g,  e�  h,  e�  n�,   "  e�	  o�,  e�  p�,  eH  v�,   *"  e`  w�,  ew  x�,  e   y�,  e~  -   5"  e   �-  e�  �-  e  �-  e�   �-  e�  �-  e�	  �-  e�  �_-   @"  e  �_-  e  �_-  e�  �_-  e�  ��-   K"  e�  ��-  e�  ��-  e�  ��-  em  ��-   V"  e	  ��-  e2	  ��-  e�  ��-  e9  ��-  e[  �
.   a"  eJ  �
.  e�  �
.  e7  �
.  e�  �?.   l"  eI	  �?.  e$	  �?.  e�   �h.   w"  eN  �h.  ep  ��.   �"  e�  ��.  e:  ��.  e�  .  ed   Å.  e�  ��.   �"  e  ��.  e�  ��.  e�	  ��.   �"  e�  ��.  e  �/   �"  e�  �/  e�  �/  e�  �/  e+  �A/   �"  e�  �A/  e�   �A/  e  �j/   �"  e�
  �j/  e�  �j/  e  �/   �"  e   �/  eF  �/  e�  �/   �"  e�  ��/  e�  ��/  eD  O�/   �"  e�  P�/  e1  Q�/  e�  W0   �"  e^  X0  e�  3+0   �"  e�  4+0  e�   8H0   #  e�  9H0  el	  =e0  #  eN  >e0  e^  ?e0  eL  @e0  ea  D�0  #  eB  E�0  e�	  F�0  e  G�0  e  H�0  ey  I�0  e�   �0   %#  e�  !�0  +�  ��  �"  1  n   g>  Y  $1  �"   h�  �1  �"    l�   � C� |� �V  C     �� (  �  �  �  E   �  �  o  �	  �  qW  !s   int   "�   �  #  .  <h   `  Ds   �  Wh   �  _z   �  es   t   ms   a  us     ~s   �  �s   3  �s   �  �s   H  �s   y  �s     �s   s  �s   T   �s   �  �s   F  �s   �  �s   �  �s     �s   V  �s   3   �  s  N:   �  V:   \	  2s   o  7s   �  <s   �  Cs   �  s   �  �  3   	pO qO !�  
std ) %@  @�  ��  Y%  !0�=  �  �b  �3   Fe  �s   �#  �  �&  �y  �3  �=  y  VB  \B   3  eq �<-  bB  �  \B  \B   lt ��1  bB  �  \B  \B   ��  eF  s   �  iB  iB  �   �K  �9  �  �  iB   �(  
!  iB    iB  �  \B   1  �A  oB  >  oB  iB  �   �5  �'  oB  b  oB  iB  �   �3  �A  oB  �  oB  �  3   +  :  3  �  uB   >  �C   �P  >  �  \B   �B  $6  bB  �  uB  uB   eof (�:  >  ?  ,N0  >  uB    E  	�  9Q  	py  G0  	sy   �T  	t�  %  	{D  J  �E   %  	�Z  e  �E  y   �:  	�b;  y  }  �  �E   �T  	�4>  �  �  �E  �   �T  	�QM  �  �  �  �E   �F  	��?  �E  �  �  �E  y    I  	�O  �E  �    �E  y   (*  	�	H      )  �E  y   �O  	�eT    A  L  �E  y   �O  	́?  y  d  o  �E  F   �$  �   �:  	Z�   _� �,   5{B  6�C  7�C  �?  �%   K  \/  E@   �e  _�  �4  c�C  �J  d�C  ��  q�  �  �C   ��  s    �C  D   W  y#  �C  s     �  �J  p�  �B  �   �   !%  �   "�B  p  �  D  �  D   #�B  �  D  s     �e  y�  $[V  �  �  !�G  !@   <  x�  �4  {�  �J  |�  �J  �A  `S  ��A  ~J  ��  �J  ��  �%  �E  �K  ��   I  ��  :!  ��C   %H  ��      %�3  2�  %�G  7�  %t3  BCD  &�'  ��O  1D  'V  ��N  bB  �  �  ND   '3  �o+  bB  �  �  ND   (�P  ��O  �  �  +D   (�M  ��P  �  �  +D   (�,  �-      +D  �   '�+  ��R  �  (  .  +D   '3  �   �  E  U  +D  D  D   �/  !�B  +D  y  �  �  D   (�O  �|6  �  �  +D  D   )(  ��6  �  �  +D  D   *�   �-  �  �  �  +D   +�1  o�*  �  �  +D  D  �    *�A  $n%  �  	  	  D   *�A  (�I  �  /	  :	  %D  �   *"A  ,�%  +D  R	  X	  D   *�1  2E)  �  p	  v	  D   *�/  6;&  �  �	  �	  D   )�>  :�>  �	  �	  %D   *S  A:2  �  �	  �	  D  �  �   )�#  K�(  �	  �	  D  �  �  �   *9  S>$  �  
  '
  D  �  �   *-U  [�7  bB  ?
  J
  D  �   ,�5  d�-  j
  �  �  �   ,	1  m�P  �
  �  �  �   ,�3  v\-  �
  �  �  3    ,nU  ��-  �
  �  �  �   ,nU  �nG  �
  �  �  �   ,nU  ��   
  �  �  �   ,nU  �IP  *  �  �  �   �J  �rR  s   I  �  �   )�=  ��H  ]  r  %D  �  �  �   )V  �)  �  �  %D   -�'  �D*  1D  .�0  ��  �  %D   /�0  ��  �  %D  D   �0  ��  �  %D  7D   �0  ��    %D  7D  �  �   �0  �  8  %D  7D  �  �  D   �0  �H  ]  %D  �  �  D   �0  �m  }  %D  �  D   �0  ��  �  %D  �  3   D   .�0  "�  �  %D  s    0�  *,Q  =D  �  �  %D  7D   0�  2�G  =D  �    %D  �   0�  =�%  =D    *  %D  3    0S� f�&  �  C  I  %D   0S� q�>  �  b  h  D   1end y<  �  �  �  %D   1end �6;  �  �  �  D   0I ��$    �  �  %D   0I ��7  �  �  �  D   0��  �lC    �    %D   0��  �CM  �    "  D   0r ��R  �  ;  A  D   0�K  �r5  �  Z  `  D   0�3  �j=  �  y    D   2�� �  �  �  %D  �  3    2�� ��F  �  �  %D  �   0I  v  �  �  �  D   2�E  �|U  �    %D  �   2�1  -�      %D   0�� 5�?  bB  7  =  D   0�:  D�6  �  V  a  D  �   0�:  UW  �  z  �  %D  �   1at k
/  �  �  �  D  �   1at ��7  �  �  �  %D  �   0�F  ��/  =D  �  �  %D  7D   0�F  �k:  =D      %D  �   0�F  ��H  =D  ,  7  %D  3    0@  DA:  =D  P  [  %D  7D   0@  U�1  =D  t  �  %D  7D  �  �   0@  )�D  =D  �  �  %D  �  �   0@  ��*  =D  �  �  %D  �   0@  �6  =D  �  �  %D  �  3    2�G  -aN      %D  3    �3  �b*  =D  7  B  %D  7D   0�3  ^ 2  =D  [  p  %D  7D  �  �   0�3  �=  =D  �  �  %D  �  �   0�3  z�T  =D  �  �  %D  �   0�3  � @  =D  �  �  %D  �  3    2� ��E  �    %D  �  �  3    0� �\+  =D  )  9  %D  �  7D   0� �u>  =D  R  l  %D  �  7D  �  �   0� g|=  =D  �  �  %D  �  �  �   0� "�@  =D  �  �  %D  �  �   0� 9k<  =D  �  �  %D  �  �  3    0� K�'  �  
    %D  �  3    0bL  d�R  =D  3  C  %D  �  �   0bL  t�2  �  \  g  %D  �   0bL  �L&  �  �  �  %D  �  �   0�%  �9F  =D  �  �  %D  �  �  7D   0�%  �|<  =D  �  �  %D  �  �  7D  �  �   0�%  ��T  =D    )  %D  �  �  �  �   0�%  ��A  =D  B  W  %D  �  �  �   0�%  b>  =D  p  �  %D  �  �  �  3    0�%  3%  =D  �  �  %D  �  �  7D   0�%  'V7  =D  �  �  %D  �  �  �  �   0�%  <�+  =D      %D  �  �  �   0�%  Q'S  =D  2  L  %D  �  �  �  3    0�%  vj.  =D  e    %D  �  �  �  �   0�%  ��9  =D  �  �  %D  �  �  �  �   0�%  �C  =D  �  �  %D  �  �  �  �   0�%  �>/  =D  �    %D  �  �  �  �   *�?  ��&  =D  0  J  %D  �  �  �  3    *�1  �O  =D  b  |  %D  �  �  �  �   ,)  �z-  �  �  �  3   D   3+E  �3J  �  �  �  3   D   0�5  ��)  �  �  �  D  �  �  �   2n	 @D      %D  =D   0W�  �6  �  *  0  D   0�A  %�A  �  I  O  D   0��  ,Z5  �  h  n  D   0�(  �;  �  �  �  D  �  �  �   0�(  I�%  �  �  �  D  7D  �   0�(  X�5  �  �  �  D  �  �   0�(  �^   �      D  3   �   0�(  v�S  �  0  @  D  7D  �   0�(  	K  �  Y  n  D  �  �  �   0�(  �o?  �  �  �  D  �  �   0�(  J5  �  �  �  D  3   �   0NW  ��Q  �  �  �  D  7D  �   0NW  /�I  �      D  �  �  �   0NW  ��,  �  0  @  D  �  �   0NW  ��;  �  Y  i  D  3   �   0�S  ��I  �  �  �  D  7D  �   0�S  >T?  �  �  �  D  �  �  �   0�S  05  �  �  �  D  �  �   0�S  $S:  �      D  3   �   0�>  2hL  �  +  ;  D  7D  �   0�>  SUB  �  T  i  D  �  �  �   0�>  Q�2  �  �  �  D  �  �   0�>  _�K  �  �  �  D  3   �   0�4  qT  �  �  �  D  7D  �   0�4  j�K  �  �    D  �  �  �   0�4  ��5  �  +  ;  D  �  �   0�4  N.  �  T  d  D  3   �   0U+  �)  4  }  �  D  �  �   0��  �!1  s   �  �  D  7D   0��  ��T  s   �  �  D  �  �  7D   0��  ��O  s   �    D  �  �  7D  �  �   0��  �;.  s   0  ;  D  �   0��  ��B  s   T  i  D  �  �  �   0��  ��,  s   �  �  D  �  �  �  �   E  !T  3   4�E  '  4�F  �   5�&  5�7  4  �o  >u"  �| Cs   6Q  b�   �  6�F c�  6�R  d�  63  e�  6�  f�  6�K  g�  6�@  h�   7all i�  ?8�� ��  !:!  ��C   !NF  ��D  !�E  ��  !p0  ��D  !�%  ��D  9S  ��D  9�R  ��D  93  ��D  9�$  ��D  9�K  ��D  9�@  ��D  9�@  ��D  )�4  �Z      TD   )�=  y)  "  (  TD   "�� 8  H  TD  �D  �   "�� X  h  TD  �  �   "�� x  �  TD  �   "N  �  �  TD  s    "�� �  �  TD  �D   )�  �U  �  �  TD  �D   *�&  �.  bB  �  �  TD   )�F  &�;  
    TD  �D  �   )�9  )�Q  .  >  TD  �D  �D   )WR  ,`2  R  b  TD  �D  �D   )�S  /=  v  �  TD  �D  �D   :e  7,  �  TD  �D  �    !�$  TD   9OD  TD  9gP  TD  9�F  $ZD  ;< �  << r�  �U  �    =id ��   !�U  ��   9�I  ��C  )�  �<?  4   ?   |D  �D   >id �N   Y   |D  �D   ?id �i   o   |D   @4H  ��(  �  �   �D    �o  u�   �   jD   �o  ~�   �   jD  pD   /�o  ��   �   jD  �   �o  ��   �   jD  pD  �  �   �o  �!  !!  jD  pD  pD  �   5  �1!  <!  jD  s    �  ��*  pD  T!  _!  jD  pD   H�  ��N  z"  w!  }!  vD   U  �9  bB  �!  �!  vD  pD   2  �t*  bB  �!  �!  vD  pD   AjP  �D  �  �!  pD   BRD  �Q  pD  C�o  7�!  
"  jD  TD   D�K  :�N  D�A  =�5  �K  @I  �  <"  �   )�,  CH<  P"  e"  jD  pD  pD  �   �  �  Q   �  � >4  EW  3#  F�4  F�$  Fq-  Fc=  Fo'  F�5   F�%  � F�8  �FX)  �F�%  �F�  �FaO  �FY=  � FP  �� F�C  ��FwS  �F�O  � F�?  �F�5  �� E
$ gM#  F)W  F�   F�U  F�A  F�8  F�P   FEH  �� E�4  �z#  FO   F�7  F(  F�Q  FG  �� E��  ��#  F�R   F�-  F�1  FlO  �� ;b4 I&  �P  ��"  G�N  �z#  G�  JM#  0n4 '�T  �#  �#  �#  �K   0�/ v2  �5  $  $  jL  �5   0l6 �6N  �5  ,$  7$  jL  �5   0-H  ��`  �  P$  V$  �K   0s0 B?  �#  o$  z$  jL  �#   0s0 S�(  �#  �$  �$  jL  �#  �#   G�9  i#  0*H  ��7  pD  �$  �$  �K   H�4  �$  �#  Idec �$  Ht-  �$  Ihex �$  Hr'  �$  H< �$   Ioct �$  @H� �$  �J[)  �$   J�%  "�$   J�  &�$   JdO  )�$   J\=  ,�$   J�P  /�$    J�C  3�$   @HzS  6�$  �H�O  9�$  JJ�?  <�$  H�7  N�%  �#  H(  Q�%  H�Q  V�%  HO  Y�%   Iin w"&  �$  Iout z"&  Icur �C&  �#   �a  $�&  rS  +a   Km�  ,l&  U&  K��  -l&  K�4  .l&  K;�  /l&  K��  0l&  K� 1l&   K�� 2l&  @Lb  3l&  L�e  4l&   L�  5l&   Kމ  6l&   �#  ;�8  ('  !T  3   4�E  '  M� �qP  �D  !'  F    N�Y  �:('  (0  8�_ ��'  !�M  �bB   G{'  �(0  Gb  ��'  GDe  �>  /�_ .�'  �'  �D  �D  bB   0�  ��e  bB  �'  �'  �D   m'  `'   b  J�2  8'  O�3  <"Pƾ �D   Q�� R�5  �b  >3   Fe  ?>  �#  @I  �&  AT  {'  E(0  �!  F�3  &� G('  F I�5  /̾ ]k(  �(  E  s   E  E   R�% g('  �(  �(  E  s   E   �� xu� E  �(  �(  E  #E   �� |׿ E  �(  �(  E  8E   �� ��� E  )  )  E  SE   �� ��� E  &)  1)  E  hE   �� �� E  I)  T)  E  nE   �� ��� E  l)  w)  E  tE   �� �ϸ E  �)  �)  E  zE   �� �K� E  �)  �)  E  �E   �� �ڸ E  �)  �)  E  �E   �� �� E  �)  *  E  �E   �� �� E  *  &*  E  �E   �� �� E  >*  I*  E  �E   �� �ĸ E  a*  l*  E  �E   �� ڮ� E  �*  �*  E  �E   �� ޹� E  �*  �*  E  �E   �� �� E  �*  �*  E  �E   0�� �� E  �*  �*  E  E   0�� �� �5  +  +  �E   1get .L� (  1+  7+  E   1get <r� E  P+  [+  E  �E   1get W�� E  t+  �+  E  �E  �5  �'   1get b3� E  �+  �+  E  �E  �5   1get yX� E  �+  �+  E  �E  �'   1get �η E  �+  �+  E  �E   0�d  j�c  �D  ,  -,  E  �E  �5  �'   0�d  �ɺ E  F,  V,  E  �E  �5   0Ic  tb  �D  o,  ,  E  �5  (   0Ic  o�d  �D  �,  �,  E  �5   0Ic  �A� E  �,  �,  E   0/� �}� (  �,  �,  E   02_  �» E  �,  
-  E  �E  �5   0� ��� �5  #-  3-  E  �E  �5   0� 
�� E  L-  W-  E  �'   0ѿ A� E  p-  v-  E   0� ,�� s   �-  �-  E   07� ;4� (  �-  �-  E   01� JӼ E  �-  �-  E  (   01� Z�� E  �-  .  E  (  �#   .̾ ^.  ".  E  s   E   O(  (  (  �� Vۺ �D  R.  ].  ]T  S   E  tE   �� Vu� �D  ~.  �.  ]T  a   E  �E   g� V�� �D  �.  �.  ]T  %   E  �E   � V�� �D  �.  �.  ]T  ,   E  �E   �� V� �D  /  /  ]T  bB  E  hE   �� V�� �D  ./  9/  ]T  �   E  �E   ߾ V� �D  Z/  e/  ]T  �   E  �E   �� VY� �D  �/  �/  ]T  <B  E  �E   j� V!� �D  �/  �/  ]T  5B  E  �E   O� V=� �D  �/  �/  ]T  .B  E  �E   � V� �D  
0  0  ]T  �  E  �E   !T  3   4�E  '   ;�M  �2  0�* �e  �F  J0  P0  �F   �b  �3   0�* �_e  �F  u0  {0  �F   0�D t> �5  �0  �0  >F   2cb  �Pc  �0  �0  >F  s    0�-  �  �F  �0  �0  �F   0�-  P  �F  �0  �0  �F   2� !4  1  1  >F  s    0% ��" �F  11  71  �F   0�a  R(b  V1  P1  V1  >F   Fe  �>  0�c  <�c  V1  {1  �1  >F   0�S  �YH  V1  �1  �1  >F  P0   0j> t�B V1  �1  �1  >F  P0   0�D �'? V1  �1  �1  >F   0�W  elD �5  2  2  >F  �F  �5   0X'  F6  s   *2  02  >F   -9  ��<  ]2  H2  ]2  >F  i2  �#  �$   �#  �I  �&  �T  0:H  ?,  ]2  �2  �2  >F  ]2  �$   0!a  *�a  V1  �2  �2  >F   !T  3   4�E  '   ;�+  t3  0��  a�)  �2  �2  �2  �L  3    G�b  �3   Sis 1�c  bB  !3  13  �L  U&  3    TKC  3�T  �2  �2  R3  ]3  �L  3    :+3  ��3  m3  �L    �� 
8�3  oS  
8�#    �� 
V�3  oS  
V�#    i� 
t�3  TC  
ts     x� 
��3  V  
�s     2� 
��3  V  
�s     ;�E  �5  03F  ;�S  >F  4  4  DF   �M  ��B  �#  14  74  DF   1tie !�G  F  P4  V4  DF   9U  ؍0  �#  n4  t4  DF   U`V  �3  �4  �4  8H  s    .aV  ��4  �4  8H   eU  ��4  �4  �4  8H  �#   0[F l�L  �4  �4  �4  DF   �b  K3   �=  �93  bB  5  5  DF   bU  �IQ  (5  35  8H  �#   Z  �4O  bB  K5  Q5  DF   0��  ��$  �4  j5  u5  DF  3    0[F ��@  �4  �5  �5  8H  �4   !T  3   4�E  '  i3 ~P4  �5  �5  8H  >F   V�1  )�%  �5  8H  �#    �>  	b�  ;�p  �8  1get �k�  26  6  26  �N  26  26  �D  HO  �E   G�B  �9  1get ��  26  X6  w6  �N  26  26  �D  HO  tE   1get ���  26  �6  �6  �N  26  26  �D  HO  �E   1get �B�  26  �6  �6  �N  26  26  �D  HO  �E   1get ���  26   7  7  �N  26  26  �D  HO  hE   1get ��  26  87  W7  �N  26  26  �D  HO  �E   1get �t�  26  p7  �7  �N  26  26  �D  HO  �E   1get y�  26  �7  �7  �N  26  26  �D  HO  �E   1get �  26  �7  �7  �N  26  26  �D  HO  �E   1get S�  26  8  78  �N  26  26  �D  HO  �E   1get 6݋  26  P8  o8  �N  26  26  �D  HO  �E   0�f  I� �A  �8  �8  |�  3   �N  �  �  3    !T  3   4�  9   ('  ��  v9  W�J  �8  �8  6N   �#    X_Tp 3   �.  �   �?  �  �   �C   ��  2�:  �8   }'  C(0  (T  a�E   Fe  B>  �>  b69  �b  @3   (� D('  X�  fv9  |9  �E   X�  p�9  �9  �E  �E   X�  t�9  �9  �E  �E   *  {p  N9  �9  �9  �E   �F  �C�  �E  �9  �9  �E   �F  �ޙ  9  :  :  �E  s    |�  ���  bB  ):  4:  �E  �E   '  �%�  69  K:  Q:  �E   '��  Ú�  bB  h:  n:  �E   69  !T  3   �E  '   9    `'  
��:  �>  
�3    !T  3    Y0T  �:  "��  :�:  �:  �W  �   !T  3    �3  (0  �5  Z�*  O�"  	;  �"  �"   Z*  K�"  #;  �"  �"   Z�*  �M#  =;  M#  M#   Z*  �M#  W;  M#  M#   Z	W  ��K  q;  �K  M#   M#  Z	W  [�K  �;  L  �"   �"  Z+  W�"  �;  �"   ZwA  _�K  �;  L  �"   �2  �  ZN  .[N  �;  �R  �2  �L   Z�� .�N  
<  �R  �5  �N   �5  Z�b  �	P  2<  X_Tp %   	P  	P   Z+  �M#  G<  M#   Z�   	�bB  j<  �$  �  F  F   ;�N  >=  0\�  �DU  z"  �<  �<  �V   0��  �  �<  �<  �<  �V   G7# p4  0�p  �kV  �<  �<  �<  �V   0�{  �w:  �<  �<  �<  �V   G�b  o3   0]�  ��H  �<  "=  (=  �V   [id >�  !T  3    j<  Z l  �bB  o=  !T  3   �E  '  �E  �E   Z��  �bB  �=  !T  3   �E  '  �E  �E   !� �l� �D  �=  !T  3   �E  '  �D   c  �� �D  �=  !T  3   �E  '  �D  �C   � ��� �D   >  �E  '  �D  �   � �Ž �D  H>  �E  '  �D  O�   � D� �D  p>  �E  '  �D  ��   � � �D  �>  �E  '  �D  �   3c  
�$� �D  �>  !T  3   �E  '  �D  �:   3c  
e�� �D  �>  !T  3   �E  '  �D  �3   3c  
G{� �D  (?  !T  3   �E  '  �D  t3   3c  
�/� �D  X?  !T  3   �E  '  �D  �3   3c  
�=� �D  �?  !T  3   �E  '  �D  �3   3c  
��� �D  �?  !T  3   �E  '  �D  �3   \	@  8�N  �U  07  �5  �?  >F  >F  hE   3}`   ��d  [N  	@  �R  �2  pD   c  da  �D  �D  �    ]$   %�.B  �  "$#,�  #-�  K  #:�A  �e  #=�  � #?�  "  #@�  �4  #A�C  �J  #B�C  �A  #O�@  �@  �C   �A  #Q�@  �@  �C  �C   �A  #V�@  �@  �C  s    �
 #Y51  ]@  �@  �@  �C  u@   �
 #]�R  i@  A  A  �C  �@   � #c?  ]@  7A  GA  �C  Q@  �   _ #m.   [A  kA  �C  ]@  Q@   �3  #q89  Q@  �A  �A  �C   .E  #��3  �A  �A  �C  ]@  �C   �(  #��(  �A  �A  �C  ]@   X_Tp 3    E@  5ZD  58E  s  $/�A  |  $0s    ^U  (A�C  B  
F  s    _9+  (N�C  
F  s     �� �� �� ]2*  !7VB  `!8    a3  ay  �  y  3  a�  �  8&�C  �{  &�   ]�  &�  \�  & �  �D  &!�  �3  &"�  U>  &#�  &�  &$�  �  &%�  �*  &&�   ڡ  &'3   $�U  &(3   %TL  &)3   &�I  &*3   'Q  &+3   (�C  &,3   )�J  &-3   *1  &.�  ,o(  &/3   0�U  &03   1PL  &13   2�I  &23   3Q  &33   4�C  &43   5�J  &53   6 Z)%  &K�  �C  s   �   bGT  &P�C  {B  �  ' s   a3   a�  E@  a�A  �A  �  a/    s   bB  @  �  4  E  aE  a�  a4  c,   ND  d �  Q  _D  eD  �  �  au"  u"  �  ae"  e"  �D  j"  �  c�D  �D  d c�D  �D  d �D  �D  ao"  o"  a�#  a�&  %   8'  a('  �'  es   �D  f E  g�5  �D  ('  �  +(  aC(  )E  eE  8E  E   >E  eME  ME  ME   a7(  YE  e�D  hE  �D   abB  aZ   aS   as   aa   a%   a,   a�   a�   a<B  a5B  a.B  a�  �8  a�'  �'  a+(  9  9  aZ9  �:  a9  a�:    �:  a  a�:  �C  h�A  >F  iXF  (A
F  i\;  (As   jk�T  (C�C    (0  �:  l�3  XF  bF  mh  bF   DF  l4  uF  F  mh  bF   �&  l74  �F  �F  mh  bF   lV4  �F  �F  mh  bF   P0  �:  l10  �F  �F  mh  �F   �F  l\0  �F  �F  mh  �F   l{0  G  G  mh  G  jn�&  �:    >F  l�0  /G  EG  mh  G  o__n �s    l�0  SG  ]G  mh  �F   l�0  kG  uG  mh  �F   l�0  �G  �G  mh  G  o__n !s    l1  �G  �G  mh  �F   hx  �G  jp__p ��    l�  �G  �G  mh  �G   D  l:	  �G  �G  mh  �G   l�  H  H  mh  H   ND  l�  )H  3H  mh  3H   +D  �3  lt4  LH  _H  mh  _H  m#  D   8H  l�(  rH  �H  mh  �H  m#  D  m�!  �H   E  E  hB  �H  iXF  (N
F  i\;  (Ns    ly  �H  �H  mh  3H  q__a ��H   D  h_  I  ihR  �I  imR  �I   VB  \B  l  I  $I  mh  3H   l�  2I  GI  mh  3H  q__n ϕ   l"  UI  _I  mh  �G   l�  mI  wI  mh  �G   h~  �I  ihR  ��I  imR  ��I   \B  \B  h�  �I  o__s 
iB  o__n 
�  o__a 
�I   \B  h�  �I  o__c �I   uB  h�  	J  o__c  	J   \B  l71  J  4J  mh  G  jn�&  TV1    lb1  BJ  ZJ  mh  G  jn�&  >V1    l�1  hJ  �J  mh  G  o__c �P0  jn�&  �V1    l�1  �J  �J  mh  G  o__c tP0  jn�&  vV1  n� wD    h�  �J  rhR  $�J  rmR  $�J   uB  uB  s�  l�1  K  #K  mh  G  jn�&  �V1    h�:  DK  q__a O�"  q__b O�"   h	;  eK  q__a K�"  q__b K�"   h#;  �K  q__a �M#  q__b �M#   h=;  �K  q__a �M#  q__b �M#   aq;  aM#  hW;  �K  q__a ��K  q__b �M#   �K  �&  l�#  �K  �K  mh  �K   �K  a�;  a�"  hv;  )L  q__a [)L  q__b [�"   L  h�;  DL  q__a W�"   h�;  eL  q__a _eL  q__b _�"   L  �#  l�#  ~L  �L  mh  �L  r�6  v�5  jn'U  x�5    jL  l$  �L  �L  mh  �L  r�R  ��5  jn'U  ��5    �;  l�2  �L  M  mh  M  o__c a3    �L  l
3  M  sM  mh  M  q__m 2U&  q__c 23   jk�&  8bB  k�`  9�;  k�b  :�  jka  =l&  jk�c  @bB      l�4  �M  �M  mh  _H   l7$  �M  �M  mh  �K   l�4  �M  �M  mh  _H  i�%  ��#   lV$  �M  �M  mh  �L  r�%  B�#  jn'U  D�#    lz$  N  6N  mh  �L  r�%  S�#  r�?  S�#  jn'U  U�#    �8  t�8  vLN  VN  mh  VN   6N  a�;  h�;  �N  �R  �2  q__f .�L   l�4  �N  �N  mh  bF   l�4  �N  �N  mh  bF   l�'  �N  �N  mh  �N   �D  a
<  
<  h�;  �N  �R  �5  q__f .�N   l�9  O  O  mh  O  q__s t�E   �E  l|9  .O  CO  mh  O  q__s pCO   �E  a�#  l�5  \O  �O  mh  �O  re  �26  r�h  �26  r$  ��O  r�*  ��O  o__v ��O   �N  �D  HO  �E  l5  �O  �O  mh  _H  i�%  ��#   l�1  �O  	P  mh  G  o__s e�F  o__n e�5   a�D  h<  9P  X_Tp %   q__a �9P  q__b �>P   	P  	P  h2<  YP  q__a �M#   l2  gP  qP  mh  G   lJ  P  �P  mh  �P  iQ  	�y   �E  l35  �P  �P  mh  bF   l02  �P  �P  mh  G  iQ  �i2  i@  ��#  i^F  ��$   l?6  �P  >Q  mh  �O  re  �26  r�h  �26  r$  �>Q  r�*  �CQ  o__v �HQ   �D  HO  tE  lw6  [Q  �Q  mh  �O  re  �26  r�h  �26  r$  ��Q  r�*  ��Q  o__v ��Q   �D  HO  �E  l�6  �Q  R  mh  �O  re  �26  r�h  �26  r$  �R  r�*  �	R  o__v �R   �D  HO  �E  l�6  !R  gR  mh  �O  re  �26  r�h  �26  r$  �gR  r�*  �lR  o__v �qR   �D  HO  hE  l7  �R  �R  mh  �O  re  �26  r�h  �26  r$  ��R  r�*  ��R  o__v ��R   �D  HO  �E  lW7  �R  -S  mh  �O  re  �26  r�h  �26  r$  �-S  r�*  �2S  o__v �7S   �D  HO  �E  l�7  JS  �S  mh  �O  re  26  r�h  26  r$  �S  r�*  �S  o__v �S   �D  HO  �E  l�7  �S  �S  mh  �O  re  26  r�h  26  r$  �S  r�*  �S  o__v �S   �D  HO  �E  l�7  T  VT  mh  �O  re  26  r�h  26  r$  VT  r�*  [T  o__v `T   �D  HO  �E  l78  sT  �T  mh  �O  re  626  r�h  626  r$  6�T  r�*  7�T  o__v 7�T   �D  HO  �E  le  �T  �T  mh  �T   �E  lu2  �T  U  mh  G  rj(  ]2  r^F  �$   hG<  ?U  �$  �  i\C  	�?U  i?)  	�DU   F  F  lo8  `U  �U  |�  3   mh  �O  �  rR'  I�  o__c I3   jn�&  Ks     �  l�  �U  �U  mh  �U  r4&  r�   �U  lQ:  �U  �U  mh  �U  jk�^  �n:    �E  l�@  �U  V  mh  V   �C  l�  V  #V  mh  #V   �C  l�@  6V  IV  mh  V  m#  D   l  WV  jV  mh  #V  m#  D   l�@  xV  �V  mh  V  �V   �C  l�  �V  �V  mh  #V  q__a s�V   D  lO  �V  �V  mh  �G   u�  �V  �V  mh  �V  m#  D   D  >=  ls<  	W  W  mh  W   �V  l�  &W  9W  mh  9W  m#  D   %D  l�<  LW  VW  mh  W   l�<  dW  nW  mh  W   l�<  |W  �W  mh  W   l	=  �W  �W  mh  W   �:  l�:  �W  �W  mh  �W  r4&  :�   �W  l`  �W  �W  mh  �V  rv�  �  o__a �W   D  s�  l�$  X   X  mh  �K   hC=  SX  !T  3   �E  '  q__a �SX  q__b �XX   �E  �E  l�9  kX  uX  mh  �U   l�9  �X  �X  mh  O   ho=  �X  !T  3   �E  '  q__a ��X  q__b ��X   �E  �E  l�  �X  �X  mh  9W   l  �X  Y  mh  9W  o__c �3    l13  Y  *Y  mh  M  o__c 33    vY  �T  ��   �EY  VY  wY  � wY  � vdH  B� ��#   �qY  �Y  xrH  lg y>H  ��   hxLH  �g z��  vdH  ��  �2   ��Y  Z  wrH  � {dH  �   h�Y  xrH  �g |>H  ��# hxLH  �g }%�  ~2���   l[(  Z  6Z  mh  �H  m#  D  m�!  6Z  i(  ]E   E  vZ  ¹ P�2   �VZ  �Z  xZ  �g x!Z  h w*Z  ����5  ���  vZ  �� ���   ��Z  [  wZ  � w*Z  �{sM  ��@   ^�Z  x�M  'h }�� {>H  �   ^�Z  wLH  s�}� ����5  � ���   vdH  A�  �   �#[  4[  wrH  � w�H  � ��(  @�   �L[  }[  �h  �H  � �$%  x#E  ��F���� �   ��(  P�   ��[  �[  �h  �H  � �$%  |8E  � ��(  p�   ��[  �[  �h  �H  � �$%  �SE  � ��*  ��   ��[  \  �h  \  �  �E  lQ5   \  6\  mh  bF  o__c �3    �-,  ��s   �N\   ]  �h  �H  � �__s ��E  ��__n ��5  ��\  ���# �]  �)\  
x \  rh �aN  ���# ��\  xtN  �h ���?   ��L  ���# �x�L  �h x�L  �h ���.   x�L  �h x�L  i ���]3     ����+   l.  .]  J]  mh  �H  m#  D  m�!  J]   E  v ]  �  �2   �j]  �]  x.]  %i x@]  9i R��5  ��0  v ]  V� `��   ��]  ^  w.]  � �sM  l�@   _�]  x�M  Mi }u� �>H  ��   _�]  wLH  s�}�� ����5  �����   l�2  ^  4^  mh  G  jn�&  ,V1    lz'   B^  �^  mh  �^  ie  /�^  i8� /bB  jk�*  1�#  jk�^  8�'  k(  9�^  p__c :m'  k�b  <�^     �D  �D  S'  �^  a�'  �4^  ѻ ���  ��^  (b  wB^  � wK^  �wV^  ��$ �b^  �i �0$ �a  �n^  �i �y^  j ��^  *j ��^  �J  v�P$ :�_  xJ  j �p$ w_  �&J  tj ��I  ��   Vx�I  �j   ���   xJ  �j ���   �&J  �j    �aN  ���$ <�_  xtN  �j ����?   �M  ���$ >�`  x*M  �k xM  l xM  Il ��$ �M  �*M  �M  ��$ �6M  4m �AM  �LM  Gm ��$ �XM  �m � % �dM  �n �K���  �����  ����  ���%�  � �:�       �^  ��@% @�a  x^  �n �@% �&^  o �4J  ��`% .6a  xBJ  �n ���   a  �LJ  Bo �!G  ��   B�/G  x8G  `o   �@�	   xBJ  to �@�	   �LJ  Bo    �J  ��x% /xJ  �o ���   �a  �&J  ��I  ��   Vx�I  �o   �p�	   xJ  �o �p�	   �&J  �o      y�I  �   ?x�I  �o   ��M  J��% Ob  x�M  1p x�M  Sp {eK  N�   �b  xzK  1p xoK  fp  ~`��5   �*�'    �1)  q��k  �Bb  fe  �h  �H  � �__n �fe  ���% Qe  ��$  v8'  �W��% Ke  ��*  y�#  �X��% �c  �__l |%   �\�ھ }ke  yp ��N  � & }�b  x�N  �p ����?   �NO  �8& ~&c  x�O  �p x�O  ]q x}O  �q �qO  �eO  x\O  yp  ��K  G�P& �oc  x�K  �q x�K  �q |eK  G�p& �xzK  �q xoK  �q   |�K  w��& �x�K  �q x�K  �q |eK  w��& �xzK  �q xoK  
r    ��M  ���& �d  x�M  r x�M  1r {eK  ��   � d  xzK  r xoK  Dr  ����5   ��& �d  ��e  ��O  ���& ��d  x�O  Xr x�O  �r {�K  ��   ��d  x�K  Xr x�K  �r yeK  ��   �xzK  Xr xoK  �r   ���O�   ���U�  ��O�  �"�i�   ��O  ��' �,e  x�O  �r x�O  s {�K  ��   �!e  x�K  �r x�K  Es yeK  ��   �xzK  �r xoK  ts   ��O�   ���U�  ��i�  �2�i�   }�� �+���  �;���   nE  pe  a".  ]  ) �e  5�  �e  a�e  �w)  �@�.  ��e  >h  �h  �H  � �__n �>h  ��0' )h  ��$  �8'  �W�X' #h  ��*  ��#  �X�x' �f  �__l �%   �\�ھ �Ch  �s ��N  u��' �Kf  x�N  �s ����?   |NO  |��' �x�O  �s x�O  Rt x}O  rt �qO  �eO  x\O  �s   ��M  ���' ��f  x�M  �t x�M  �t {eK  ��   ��f  xzK  �t xoK  �t  ����5   ��' �g  �Hh  ��O  � ( �lg  x�O  �t x�O  �t {�K  �   �ag  x�K  �t x�K   u yeK  �   �xzK  �t xoK  Ou   ��O�   ��U�  �K�O�  �U�i�   ��O  &�( �h  x�O  cu x�O  �u {�K  .�   ��g  x�K  cu x�K  �u yeK  .�   �xzK  cu xoK  �u   �P�O�   �$�U�  �=�i�  �e�i�   }X� �^���  �n���   zE  pe  �e  ��*  �p�  �gh  |j  �h  �H  � ��D  E  ��8( gj  ��*  ��#  �u ��$  �8'  �n�X( �h  �Z*  �bB  �o����?   �p( yi  �|j  ��O  ��( �Zi  x�O  3v x�O  _v {�K  �   �Oi  x�K  3v x�K  �v yeK  �   �xzK  3v xoK  �v   �#�O�   ��U�  �P�O�  �Z�i�   ��O  .��( ��i  x�O  �v x�O  �v {�K  6�   ��i  x�K  �v x�K  w yeK  6�   �xzK  �v xoK  7w   �U�O�   ��M  ���( �Cj  ��M  x�M  Kw {eK  ��   �8j  �zK  xoK  ^w  ����5   }���,�U�  �E�i�  �j�i�   �c���  �s���   �e  �+  ��0  ��j  8m  �h  �H  � ��( #m  ��^  �'.  �__c �(  rw ��*  ��#  �w ��$  �8'  �o�4J  ��) ��k  xBJ  �w ���   dk  �LJ  �w ��I  ��   ABk  x�I  x  �!G  ��   B�/G  x8G  4x   �0�   xBJ  Hx �0�   �LJ     ��O  �� ) l  x�O  [x x�O  �x {�K  ��   ��k  x�K  [x x�K  �x yeK  ��   �xzK  [x xoK  �x   ���O�   �@) �l  �8m  ��O  o�X)  �l  x�O  �x x�O  �x {�K  u�   ��l  x�K  �x x�K  y yeK  u�   �xzK  �x xoK  ;y   ���O�   �m�U�  ���O�  ���i�   ��M  �p) 	�l  ��M  x�M  Oy {eK  �   ��l  �zK  xoK  by  ���5   }�����U�  ���i�  ���i�   �����  �����   �e  �7+  ��  �Xm  !p  �h  �H  � �__c <!p  ���) p  ��*  �#  vy ��$  8'  �o� �A   sn  n�1 '.  �4J  ��) Wn  xBJ  �y ��   1n  �LJ  �y ��I  �   An  x�I  �y  �!G  �   B�/G  x8G  	z   �0�   xBJ  z �0�   �LJ     ��I  ��) x�I  0z   ��) o  �&p  ��O  _��) %�n  x�O  Hz x�O  tz {�K  e�   ��n  x�K  Hz x�K  �z yeK  e�   �xzK  Hz xoK  �z   �t�O�   �]�U�  ���O�  ���i�   ��O  �* )�o  x�O  �z x�O  { {�K  ��   ��o  x�K  �z x�K  *{ yeK  ��   �xzK  �z xoK  L{   ���O�   ��M  ��0* .�o  ��M  x�M  `{ {eK  ��   ��o  �zK  xoK  s{  ����5   }���}�U�  ���i�  ���i�   �����  �����   �E  �e  �[+  4���  �Fp  �t  �h  �H  � �__s W�E  �{ �__n W�5  ���e  W�'  ��H* ot  ��*  8�#  �{ ��$  98'  �_�h* �r  ��a  >'.  :| ��^  ?'.  q| �(  @E  �| �__c A(  �| ��I  �   >q  x�I  �|  �J  �   ALq  xJ  �| ��   �&J    �^   ��* Ijr  x^  7} ��* �&^  `} �J   ��* /�q  xJ  �} � �   �q  xJ  �} � �   �&J    �e�   �&J  ��I  i�   Vx�I  �}    �4J  [��* .xBJ  7} �[�
   Br  �LJ  �} �!G  _�   B�/G  x8G  �}   ���   xBJ  �} ���   �LJ       ��I  N�	   G�r  x�I  ~  ��K  |�   L��K  ��K    ��* Qs  ��t  ��O  ��* P2s  x�O  P~ x�O  |~ {�K  !�   �'s  x�K  P~ x�K  �~ yeK  !�   �xzK  P~ xoK  �~   �0�O�   ��U�  �b�O�  �l�i�   ��O  ;�+ T�s  x�O  �~ x�O   {�K  C�   ��s  x�K  �~ x�K  = yeK  C�   �xzK  �~ xoK  l   �g�O�   ��K  ��   [�s  x�K  � x�K  �  ��M  ��(+ ]Kt  x�M  � x�M  � {eK  ��   �@t  xzK  � xoK  �  ����5   }���9�U�  �R�i�  �|�i�   �u���  �����   �e  ��+  ��s   ��t  su  �h  �H  � �__s b�E  ��__n b�5  ��\  ��@+ chu  �)\  
x \  � �aN  ��X+ �u  xtN  "� ���?   ��L  ��p+ �x�L  @� x�L  T� ���.   x�L  r� x�L  �� ���]3     ���+p   ��+  c�
  ��u  Lz  �h  �H  � �(  yLz  ���e  y�'  ���+ 7z  ��*  g�#  �� ��$  h8'  �_��+ �x  ��a  m'.  р ��^  n'.  � �`� oE  @� �__c p(  t� �mR  q�'  �� ��I  ?�   mdv  x�I  �  �J  S��+ p�v  xJ  @� �S�   �v  �&J  L� ��I  \�   Vx�I  j�   ��+ xJ  }� ��+ �&J     ��I  g�   q�v  x�I  ��  �ZJ  v��+ u�w  xqJ  Ȃ xhJ  � �v�   Tw  �~J  � �uG  ��
   ���G  x�G  $�   �p�   xqJ  8� xhJ  K� �p�   �~J  ��I  v�   �x�I  j�     �^  ���+ xx^  �� ��+ �&^  �� �4J  ��, .Fx  xBJ  �� ���    x  �LJ  ̓ �!G  ��   B�/G  x8G  ��   � �   xBJ  � � �   �LJ     �J  ��(, /xJ  � ���   ux  �&J   �@�0   xJ  %� �@�0   �&J        ��O  ��@, �y  x�O  8� x�O  d� {�K  ��   �y  x�K  8� x�K  �� yeK  ��   �xzK  8� xoK  ��   ���O�   �`, �y  �Qz  ��O  ��x, ��y  x�O  Є x�O  �� {�K  ��   ��y  x�K  Є x�K  � yeK  ��   �xzK  Є xoK  0�   ���O�   ���U�  ���O�  ��i�   ��M  ���, �z  ��M  x�M  D� {eK  �   �z  �zK  xoK  W�  ���5   }2����U�  ���i�  ��i�   �
���  ����   �E  �e  ��+   �s   �nz  0{  �h  �H  � �(  �0{  ��\  +��, �%{  �)\  
x \  k� �aN  2��, ��z  xtN  �� ����?   ��L  6��, �x�L  Ņ x�L  م �`�.   x�L  �� x�L  � �i�]3     �N�su   �E  ��,  ���  �P{  �}  �h  �H  � ��, �}  ��$  �8'  �o�- �}  ��*  ��#  � �0- 6|  ��^  �'.  �(  �E  J� �4J  ��H- �xBJ  J� ���   |  �LJ  h� �!G  ��   B�/G  x8G  {�   � �   xBJ  �� � �   �LJ      ��M  �`- ��|  x�M  �� x�M  �� {eK  �   ��|  xzK  �� xoK  Ɇ  �(��5   �x- 7}  ��}  ��O  =��- �}  x�O  ݆ x�O  	� {�K  C�   �}  x�K  ݆ x�K  2� yeK  C�   �xzK  ݆ xoK  a�   �R�O�   �;�U�  ���O�  ���i�   ��O  ]��- ��}  x�O  u� x�O  �� {�K  e�   ��}  x�K  u� x�K  �� yeK  e�   �xzK  u� xoK  �   ���O�   �[�U�  �t�i�  ���i�   }�� �����  �����   �e  ��,  k���   �~  ��  �h  �H  � ��- v�  �__c n(  �� ��$  p8'  �o��- p�  ��*  s�#  G� �J  �� . v�~  xJ  �� ���   �~  �&J  �� ��I  ��   Vx�I  Ԉ   ���   xJ  � ���   �&J     ��M  �8. �.  x�M  �� x�M  � {eK  �   �#  xzK  �� xoK  !�  ���5   ��O  /�P. ��  x�O  5� x�O  a� {�K  5�   ��  x�K  5� x�K  �� yeK  5�   �xzK  5� xoK  ��   ���O�   �p. Q�  ���  ��O  g��. |2�  x�O  ͉ x�O  � {�K  m�   �'�  x�K  ͉ x�K  � yeK  m�   �xzK  ͉ xoK  -�   �|�O�   �e�U�  ���O�  ���i�   �-�U�  �D�i�  ���i�   }�� �����  �����   �e  ��,  ����   ���  �  �h  �H  � �__s ��E  ��__n ��5  ���. ނ  ��$  �8'  �o��. ؂  ��*  ��#  A� ��O  ��   �>�  x�O  m� x�O  �� x�O  Ŋ  ��M  ��. ���  x�M  ؊ x�M  � {eK  �   ���  xzK  ؊ xoK  ��  ���5   �/ ?�  ��  ��O  4�0/ � �  x�O  � x�O  ?� {�K  :�   ��  x�K  � x�K  h� yeK  :�   �xzK  � xoK  ��   �I�O�   �2�U�  �y�O�  ���i�   ��O  T�H/ ���  x�O  �� x�O  ׋ {�K  \�   ���  x�K  �� x�K  �� yeK  \�   �xzK  �� xoK  �   �~�O�   �R�U�  �k�i�  ���i�   }�� �����  �����   �e  �
-  ���:  ��  ͅ  �h  �H  � �__s ��E  ��__n ��5  ��h/ ��  ��$  �8'  �o��/ ��  ��*  ��#  +� ��/ �  �	e  ��:  c� ��F  ���/ ��  xG  �� ���
   ǃ  �G  ��  � �   xG  ڌ � �   �G     ��O  ���/ ���O  x�O  � x�O  �   ��M  B� 0 �p�  x�M  ,� x�M  @� {eK  J�   �e�  xzK  ,� xoK  S�  �W��5   �0 �  �ͅ  ��O  o�80 ���  x�O  g� x�O  �� {�K  u�   ��  x�K  g� x�K  �� yeK  u�   �xzK  g� xoK  �   ���O�   �m�U�  ���O�  ���i�   ��O  ��P0 ���  x�O  �� x�O  +� {�K  ��   ���  x�K  �� x�K  I� yeK  ��   �xzK  �� xoK  k�   ���O�   ���U�  ���i�  ���i�   }�� �����  �����   �e  �3-  ���  ��  �  �h  �H  � �__c 
�'  ��p0 ��  ��$  �8'  �o��K  ��   �J�  ��K  }x�K  �  ��0 ��  ��*  ��#  �� ��0 E�  ��^  �'.  �� �(  �E  Վ ��J  2��0 �x�J  � x�J  2� ��0 �  ��J  P� ��J  c� �!G  ��   }�/G  x8G  �   �>�   x�J  �� x�J  3� �>�   ��J  ��J  ��I  @��0 zx�I  F�      ��M  `�   ���  x�M  n� x�M  �� �eK  `� 1 ���  xzK  n� xoK  ��  �p��5   �1 G�  ��  ��O  ��81 �(�  x�O  �� x�O  Ր {�K  ��   ��  x�K  �� x�K  �� yeK  ��   �xzK  �� xoK  -�   ���O�   ���U�  ���O�  ���i�   ��O  ��P1 ���  x�O  A� x�O  m� {�K  ��   ���  x�K  A� x�K  �� yeK  ��   �xzK  A� xoK  ��   ���O�   ���U�  ���i�  ���i�   �	��5  }� �����  �����   �e  �W-  � �  �%�  �  �h  �H  � �p1 ߋ  ��$  �8'  �o��K  �   �r�  ��K  }x�K  ��  ��1 ϋ  ��*  ��#  Ց ��1 4�  ��^  �'.  � �(  �E  #� ��J  N��1 �xK  A� �N�   �  �K  _� �!G  S�   ��/G  x8G  r�   �`�   xK  �� �`�   �K      ��M  ���1 ��  x�M  �� x�M  �� �eK  ��2 ���  xzK  �� xoK  ��  ����5   � 2 6�  ��  ��O  ��@2 ��  x�O  Ւ x�O  � {�K  ��   ��  x�K  Ւ x�K  *� yeK  ��   �xzK  Ւ xoK  Y�   ���O�   ���U�  ���O�  ���i�   ��O  ��X2 ��  x�O  m� x�O  �� {�K  ��   ���  x�K  m� x�K  �� yeK  ��   �xzK  m� xoK  ٓ   ���O�   ���U�  ���i�  �	�i�   �%��5  }4� ����  ����   �e  �v-   ��   ��  W�  �h  �H  � �x2 B�  ��&  s   � ��$  8'  �o��2 <�  ��*  �#  � �?�    ��  �(  E  R� �YP  L�   xgP  e�   ��M  ���2 )��  x�M  x� x�M  �� {eK  ��   ��  xzK  x� xoK  ��  ����5   ��2 ��  �W�  ��O  ��3 #��  x�O  �� x�O  ߔ {�K  ��   �y�  x�K  �� x�K  � yeK  ��   �xzK  �� xoK  7�   ���O�   ���U�  ���O�  ��i�   ��O  �� 3 '�  x�O  K� x�O  w� {�K  ��   ��  x�K  K� x�K  �� yeK  ��   �xzK  K� xoK  ϕ   ���O�   ���U�  ���i�  ��i�   }6� ����  ����   �e  ��-  0 ��   �w�  e�  �h  �H  ��@3 P�  ��&  5(  � ��$  68'  �c�qP  1�   5Վ  ��P  xP  �  ��P  s�h3 <	�  ��P  ��P  ��P   x�P  v�  ��3 ��  �e�  ��O  ���3 A��  x�O  �� x�O  �� {�K  ��   ���  x�K  �� x�K  ޖ yeK  ��   �xzK  �� xoK  �   ���O�   ���U�  ���O�  ��i�   ��O  ���3 E,�  x�O  !� x�O  M� {�K  ��   �!�  x�K  !� x�K  v� yeK  ��   �xzK  !� xoK  ��   � �O�   }G����U�  ���i�  ��i�   ����  ����   �e  ��-  L �  ���  �  �h  �H  � �%  J(  ���3 �  ��$  S8'  �G��K  3�   R�  ��K  }x�K  ��  ��3 ��  ��*  V�#  ͗ �v�/   F�  �__p \,.  �H��T  v�4 ]�U  w�T  �Tx�T  �   ��M  �� 4 l��  x�M  0� x�M  D� {eK  ��   ���  xzK  0� xoK  W�  ����5   �84 G�  ��  ��O  ��X4 f(�  x�O  k� x�O  �� {�K  ��   ��  x�K  k� x�K  �� yeK  ��   �xzK  k� xoK  �   ���O�   ���U�  ��O�  � �i�   ��O  ��p4 j��  x�O  � x�O  /� {�K  ��   ���  x�K  � x�K  M� yeK  ��   �xzK  � xoK  o�   ��O�   ���U�  ��i�  �0�i�   �@��5  }O� �)���  �9���   �e  ��-  s@�  �%�  ��  �h  �H  � �Q  Z(  ���J  Z�#  ���4 ��  ��$  z8'  �S��K  Y�   y��  ��K  }x�K  ��  ��4 ��  ��*  }�#  �� ���"   �  �__p �,.  �T��P  ���4 ���P  w�P  uw�P  V�W�x�P  ϙ   ��M  ���4 �Z�  x�M  � x�M  �� {eK  ��   �O�  xzK  � xoK  	�  ����5   ��4 �  ���  ��O  ��5 ��  x�O  � x�O  I� {�K  ��   �ٔ  x�K  � x�K  r� yeK  ��   �xzK  � xoK  ��   ��O�   ���U�  �6�O�  �@�i�   ��O  �(5 �}�  x�O  �� x�O  � {�K  �   �r�  x�K  �� x�K  
� yeK  �   �xzK  �� xoK  9�   �;�O�   ��U�  �(�i�  �P�i�   �f��5  }u� �I���  �Y���   �e  v�N  �e  `�   ��  �  w�N  �  ��=  p�W  ���  !T  3   �E  '  �e  ���  � �H5 ��  �{'  �(0  �De  �(  �b  ��2  ��b  �b�  M� g�  am�  D�  ��^   ��  x� 7�  �(  ��  �� *�  �__c 7�  � ��M  v�x5 �Ԗ  x�M  &� }�� �J  ���5 H�  xJ  �� ��5 �  �&J  ��I  ��   Vx�I  D�   �� 	   xJ  W� �� 	   �&J  j�    �M  ���5 �  x*M  }� xM  �� xM  ֜ ��5 �M  �*M  �M  ��5 �6M  
� �AM  �LM  � �6 �XM  �� �86 �dM  ^� �y���  �����  ����  ���%�  � :�       �^  	�X6 )�  x^  �� �X6 �&^  � �4J  	��6 .��  xBJ  �� �	�   ��  �LJ  '� �!G  �	   B�/G  x8G  E�   �0    xBJ  Y� �0    �LJ  '�    �J  ��6 /xJ  y� ��6 ��  �&J  ��I  %�   Vx�I  ��   �p    xJ  �� �p    �&J  ��      ��I  /�   H�  x�I  ӟ  ��M  J �6 	��  x�M  � x�M  � {eK  R    ���  xzK  � xoK  2�  �_ �5   ����?  }��}�  �� ��   �D  ��=  �   �֜  !T  3   �E  '  �e  �֜  � �__c �ۜ  ���6 ��  �De  �(  ��$  �8'  �o�7 ��  ��*  ��#  F� �07 !�  n�1 �c�  �  �4J  H7 ��  xBJ  r� �   ߚ  �LJ  �� ��I     A��  x�I  ��  �!G     B�/G  x8G  ͠   �0   xBJ  � �0   �LJ     ��I     �x�I  ��   ��M  C`7 �y�  x�M  � x�M   � {eK  K   �n�  xzK  � xoK  3�  �X�5   �x7 "�  ���  ��O  m�7 ��  x�O  G� x�O  s� {�K  s   ���  x�K  G� x�K  �� yeK  s   �xzK  G� xoK  ˡ   ��O�   �kU�  ��O�  ��i�   ��O  ��7 ���  x�O  ߡ x�O  � {�K  �   ���  x�K  ߡ x�K  )� yeK  �   �xzK  ߡ xoK  K�   ��O�   ��U�  ��i�  ��i�   }�  ����  ����   �D  �C  �e  aE   ��=  �   �E�  �E  '  �e  �E�  � �__c �J�  ��ř  �� � ���  �D  �  aL   � >  �   ���  �E  '  �e  ���  � �__c ���  ��ř  �� � ���  �D  O�  E   �H>      ��  �E  '  �e  �  � �__s ��  �	@  �� � ���  �D  L   �p>     �~�  �E  '  �e  ~�  � �__s �  �	@  �� � ���  �D  lu5  ��  ��  mh  _H  r�R  ��4  jn'U  ��4    ��>   z   �ߟ  !T  3   �E  '  �]\  
�ߟ  _� �__f 
��:  �� |��  .�7 
�w��  �x��  ע ��7 ���   � ��N  .�7 �x�N  ע �\  P8 p�)\   x \  "� �aN  S08 ���  xtN  @� ���?   ��L  WH8 �x�L  ^� x�L  s� �p%   x�L  �� x�L  �� �y]3         �D  ��>  �   ���  !T  3   �E  '  �]\  
e��  � �__f 
e�3  �� y�M  �   
gw�M  �w�M  R��   ��M  أ �L  �   EwL  �wL  r�y#K  �   \w8K  �x-K  أ      �D  ��>  �   ���  !T  3   �E  '  �]\  
G��  � �__f 
Gt3  �|�M  �`8 
IxN  � �N   wN  Q�`8 �(N  � �.L  �x8 V@�  x8L  �  �DL  �   VxYL  � wNL  q�yDK  �   `xYK  � xNK  �      �D  �(?  �G   ���  !T  3   �E  '  �]\  
���  @� �__f 
��3  _� y�M  
   
�xN  �� �N  xN  �� �
   �(N  Ǥ �DL  
   VY�  xYL  ۤ xNL  � yDK  
   `xYK  ۤ xNK  Ǥ   �L     WxL  � xL  � y#K     \x8K  � x-K  0�      �D  �X?  0   ��  !T  3   �E  '  �]\  
��  � �__f 
ȿ3  e� |pL  4�8 
�x~L  �� w�L  ���8 ��L  ��    �D  ��?  P   ���  !T  3   �E  '  �]\  
朣  � �__f 
��3  ҥ |�L  T�8 
�x�L  � w�L  ���8 ��L   �    �D  �1.  p  �£  H�  ]T  S   �h  �H  � �__v WH�  ���8 3�  ��$  Y8'  �[��8 -�  ��*  \�#  �\�9 ��  �ھ _M�  ?� ��N  �(9 _R�  x�N  R� ��?   y�P  �,   `x1Q  p� x%Q  �� xQ  � �Q  xQ  x� x�P  ?�   ��M  �@9 j�  x�M  Ч x�M  � {eK  �   ��  xzK  Ч xoK  �  ��5   �X9 ��  �R�  ��O  &x9 dv�  x�O  � x�O  B� {�K  ,   �k�  x�K  � x�K  k� yeK  ,   �xzK  � xoK  ��   �;O�   �$U�  �kO�  �ui�   ��O  F�9 h�  x�O  �� x�O  ڨ {�K  N   ��  x�K  �� x�K  � yeK  N   �xzK  �� xoK  2�   �pO�   �DU�  �]i�  ��i�   }� �~��  ����   tE  pe  �e  �T)  �   �o�  ��  �h  �H  � �__n ���  ����  �� � ���  tE  �].  �  �Φ  T�  ]T  a   �h  �H  � �__v WT�  ���9 ?�  ��$  Y8'  �[��9 9�  ��*  \�#  �\��9 ��  �ھ _Y�  F� ��N  �: _^�  x�N  Y� �F�?   yMQ  �,   `x�Q  w� x�Q  �� x|Q  � �pQ  xdQ  � x[Q  F�   ��M  "0: j��  x�M  ת x�M  �� {eK  *   ��  xzK  ת xoK  	�  �4�5   �H: ��  �^�  ��O  Vh: d��  x�O  � x�O  I� {�K  \   �w�  x�K  � x�K  r� yeK  \   �xzK  � xoK  ��   �kO�   �TU�  ��O�  ��i�   ��O  v�: h�  x�O  �� x�O  � {�K  ~   ��  x�K  �� x�K  
� yeK  ~   �xzK  �� xoK  9�   ��O�   �tU�  ��i�  ��i�   }� ����  ����   �E  pe  �e  ��)  �   �{�  ��  �h  �H  � �__n ���  ����  �� � ���  �E  ��.  �  �ک  `�  ]T  %   �h  �H  � �__v W`�  ���: K�  ��$  Y8'  �[��: E�  ��*  \�#  �\��: ��  �ھ _e�  M� ��N  ; _j�  x�N  `� �v�?   yNO  ,   `x�O  ~� x�O  �� x}O  � �qO  xeO  �� x\O  M�   ��M  R ; j�  x�M  ޭ x�M  �� {eK  Z   ���  xzK  ޭ xoK  �  �d�5   �8; ��  �j�  ��O  �X; d��  x�O  $� x�O  P� {�K  �   ���  x�K  $� x�K  y� yeK  �   �xzK  $� xoK  ��   ��O�   ��U�  ��O�  ��i�   ��O  �p; h&�  x�O  �� x�O  � {�K  �   ��  x�K  �� x�K  � yeK  �   �xzK  �� xoK  @�   ��O�   ��U�  ��i�  ��i�   }� ����  ����   �E  pe  �e  ��)  �   ���  ��  �h  �H  � �__n ���  ����  �� � ���  �E  ��.     ��  l�  ]T  ,   �h  �H  � �__v Wl�  ���; W�  ��$  Y8'  �[��; Q�  ��*  \�#  �\��; ��  �ھ _q�  T� ��N  7�; _v�  x�N  g� ���?   y�Q  ;,   `x�Q  �� x�Q  �� x�Q  &� ��Q  x�Q  �� x�Q  T�   ��M  �< j�  x�M  � x�M  � {eK  �   ��  xzK  � xoK  �  ���5   �(< ��  �v�  ��O  �H< d��  x�O  +� x�O  W� {�K  �   ���  x�K  +� x�K  �� yeK  �   �xzK  +� xoK  ��   ��O�   ��U�  ��O�  �i�   ��O  �`< h2�  x�O  ñ x�O  � {�K  �   �'�  x�K  ñ x�K  � yeK  �   �xzK  ñ xoK  G�   � O�   ��U�  ��i�  �i�   } ���  ���   �E  pe  �e  ��)      ���  ̯  �h  �H  � �__n �̯  �%Ŭ  �� � ���  �E  ��.  0  ��  x�  ]T  bB  �h  �H  � �__v Wx�  ���< c�  ��$  Y8'  �[��< ]�  ��*  \�#  �\��< ư  �ھ _}�  [� ��N  g�< _��  x�N  n� ���?   yR  k,   `xZR  �� xNR  �� xBR  -� �6R  x*R  �� x!R  [�   ��M  � = j�  x�M  � x�M  � {eK  �   ��  xzK  � xoK  �  ���5   �= ű  ���  ��O  �8= d��  x�O  2� x�O  ^� {�K  �   ���  x�K  2� x�K  �� yeK  �   �xzK  2� xoK  ��   ��O�   ��U�  �+	O�  �5	i�   ��O  	P= h>�  x�O  ʴ x�O  �� {�K  	   �3�  x�K  ʴ x�K  � yeK  	   �xzK  ʴ xoK  N�   �0	O�   �	U�  �	i�  �E	i�   }H �>	��  �N	��   hE  pe  �e  �)  P	   ���  ز  �h  �H  � �__n �ز  �U	ѯ  �� � ���  hE  �/  `	  ���  ��  ]T  �   �h  �H  � �__v W��  ��p= o�  ��$  Y8'  �[��= i�  ��*  \�#  �\��= ҳ  �ھ _��  b� ��N  �	�= _��  x�N  u� �
�?   yvR  �	,   `x�R  �� x�R  �� x�R  4� ��R  x�R  �� x�R  b�   ��M  �	�= j)�  x�M  � x�M  � {eK  �	   ��  xzK  � xoK  %�  ��	�5   �> Ѵ  ���  ��O  
(> d��  x�O  9� x�O  e� {�K  
   ���  x�K  9� x�K  �� yeK  
   �xzK  9� xoK  ��   �+
O�   �
U�  �[
O�  �e
i�   ��O  6
@> hJ�  x�O  ѷ x�O  �� {�K  >
   �?�  x�K  ѷ x�K  &� yeK  >
   �xzK  ѷ xoK  U�   �`
O�   �4
U�  �M
i�  �u
i�   }x	 �n
��  �~
��   �E  pe  �e  �*  �
   ���  �  �h  �H  � �__n ��  ��
ݲ  �� � ���  �E  �9/  �
  �
�  ��  ]T  �   �h  �H  � �__v W��  ��`> {�  ��$  Y8'  �[��> u�  ��*  \�#  �\��> ޶  �ھ _��  i� ��N  �
�> _��  x�N  |� �6�?   y�R  �
,   `x S  �� xS  �� xS  ;� ��R  x�R  �� x�R  i�   ��M  �> j5�  x�M  �� x�M  � {eK     �*�  xzK  �� xoK  ,�  �$�5   ��> ݷ  ���  ��O  F? d��  x�O  @� x�O  l� {�K  L   ���  x�K  @� x�K  �� yeK  L   �xzK  @� xoK  ĺ   �[O�   �DU�  ��O�  ��i�   ��O  f0? hV�  x�O  غ x�O  � {�K  n   �K�  x�K  غ x�K  -� yeK  n   �xzK  غ xoK  \�   ��O�   �dU�  �}i�  ��i�   }�
 ����  ����   �E  pe  �e  �&*  �   ���  �  �h  �H  � �__n ��  ���  �� � ���  �E  �e/  �  ��  ��  ]T  <B  �h  �H  � �__v W��  ��P? ��  ��$  Y8'  �[�x? ��  ��*  \�#  �\��? �  �ھ _��  p� ��N  ��? _��  x�N  �� �f�?   y<S  �,   `x�S  �� xwS  �� xkS  B� �_S  xSS  �� xJS  p�   ��M  B�? jA�  x�M  � x�M   � {eK  J   �6�  xzK  � xoK  3�  �T�5   ��? �  ���  ��O  v@ dʺ  x�O  G� x�O  s� {�K  |   ���  x�K  G� x�K  �� yeK  |   �xzK  G� xoK  ˽   ��O�   �tU�  ��O�  ��i�   ��O  � @ hb�  x�O  ߽ x�O  � {�K  �   �W�  x�K  ߽ x�K  4� yeK  �   �xzK  ߽ xoK  c�   ��O�   ��U�  ��i�  ��i�   }� ����  ����   �E  pe  �e  �I*  �   �û  ��  �h  �H  � �__f ���  ����  �� � ���  �E  ��/  �  �"�  ��  ]T  5B  �h  �H  � �__v W��  ��@@ ��  ��$  Y8'  �[�h@ ��  ��*  \�#  �\��@ ��  �ھ _��  w� ��N  '�@ _��  x�N  �� ���?   y�S  +,   `x�S  �� x�S  �� x�S  I� ��S  x�S  �� x�S  w�   ��M  r�@ jM�  x�M  � x�M  '� {eK  z   �B�  xzK  � xoK  :�  ���5   ��@ ��  ���  ��O  ��@ dֽ  x�O  N� x�O  z� {�K  �   �˽  x�K  N� x�K  �� yeK  �   �xzK  N� xoK  ��   ��O�   ��U�  ��O�  ��i�   ��O  �A hn�  x�O  �� x�O  � {�K  �   �c�  x�K  �� x�K  ;� yeK  �   �xzK  �� xoK  j�   ��O�   ��U�  ��i�  �i�   } ����  ���   �E  pe  �e  �l*     �Ͼ  �  �h  �H  � �__f ��  ��  �� � ���  �E  ��/     �.�  ��  ]T  .B  �h  �H  � �__v W��  ��0A ��  ��$  Y8'  �[�XA ��  ��*  \�#  �\�xA �  �ھ _��  ~� ��N  W�A _��  x�N  �� ���?   yT  [,   `xIT  �� x=T  �� x1T  P� �%T  xT  �� xT  ~�   ��M  ��A jY�  x�M  � x�M  .� {eK  �   �N�  xzK  � xoK  A�  ���5   ��A �  ���  ��O  ��A d��  x�O  U� x�O  �� {�K  �   ���  x�K  U� x�K  �� yeK  �   �xzK  U� xoK  ��   ��O�   ��U�  �O�  �%i�   ��O  � B hz�  x�O  �� x�O  � {�K  �   �o�  x�K  �� x�K  B� yeK  �   �xzK  �� xoK  q�   � O�   ��U�  �i�  �5i�   }8 �.��  �>��   �E  pe  �e  ��*  @   ���  �  �h  �H  � �__f ��  �E�  �� � ���  �E  ��/  P  �:�  ��  ]T  �  �h  �H  � �__v W��  �� B ��  ��$  Y8'  �[�HB ��  ��*  \�#  �\�hB �  �ھ _��  �� ��N  ��B _��  x�N  �� ���?   yeT  �,   `x�T  �� x�T  �� x�T  W� ��T  x|T  �� xsT  ��   ��M  ��B je�  x�M  � x�M  5� {eK  �   �Z�  xzK  � xoK  H�  ���5   ��B �  ���  ��O  �B d��  x�O  \� x�O  �� {�K     ���  x�K  \� x�K  �� yeK     �xzK  \� xoK  ��   �O�   �U�  �KO�  �Ui�   ��O  &�B h��  x�O  �� x�O   � {�K  .   �{�  x�K  �� x�K  I� yeK  .   �xzK  �� xoK  x�   �PO�   �$U�  �=i�  �ei�   }h �^��  �n��   �E  pe  �e  ��*  p   ���   �  �h  �H  � �__p � �  �u�  �� � ���  �E  �U  =2�   �   ��   >2�  �B  ?2�  ��  E^�   �   �B   F^�  �C  G^�  �e  H^�  �8  I^�  ��  J^�  �

  X��   �   ��  Y��  ��
  Z��  ��   `��  �   ��  f��   �   ��  g��  ��  h��  ��  n�   �   ��	  o�  ��  p�  �H  vG�   �   �`  wG�  �w  xG�  �   yG�  �~  ��   �   �   ���  ��  ���  �  ���  ��   ���  ��  ���  ��	  ���  ��  ���   �   �  ���  �  ���  ��  ���  ��  ��   �   ��  ��  ��  ��  ��  ��  �m  �R�     �	  �R�  �2	  �R�  ��  �R�  �9  �R�  �[  ���     �J  ���  ��  ���  �7  ���  ��  ���     �I	  ���  �$	  ���  ��   ���   "  �N  ���  �p  ��   -  ��  ��  �:  ��  ��  ��  �d   ��  ��  �b�   8  �  �b�  ��  �b�  ��	  ю�   C  ��  Ҏ�  �  ح�   N  ��  ٭�  ��  ڭ�  ��  ۭ�  �+  ���   Y  ��  ���  ��   ���  �  ��   d  ��
  ��  ��  ��  �  �>�   o  �   �>�  �F  �>�  ��  �j�   z  ��  �j�  ��  �j�  �D  O��   �  ��  P��  �1  Q��  ��  W��   �  �^  X��  ��  3��   �  ��  4��  ��   8 �   �  ��  9 �  �l	  =�  �  �N  >�  �^  ?�  �L  @�  �a  DX�  �  �B  EX�  ��	  FX�  �  GX�  �  HX�  �y  IX�  ��   ��   �  ��  !��  �  *�1  ��  �   �>  Y  ��  �   Z�e  +rs   ��  s    Zb  +^s   �  s    Z�e  +Js   %�  s    ZWe  +|s   :�  s    Z�d  +�s   O�  s    ��  ��  �  i�  �   ��   �2   �# K� � �V  HE     p� (  _� �7   �  �  �  P   �  �  o  �	  �  qW  !~   int   "�   �  #  .  <s   `  D~   �  Ws   �  _�   �  e~   t   m~   a  u~     ~~   �  �~   3  �~   �  �~   H  �~   y  �~     �~   s  �~   T   �~   �  �~   F  �~   �  �~   �  �~     �~   V  �~   >   �  s  NE   �  VE   \	  2~   o  7~   �  <~   �  C~   �  ~   �  �  >   pO qO !�  	std  c$  
@  %  0�=  	��  �b  	�>   Fe  	�~   �3  	�=  d  k(  q(   4  eq 	�<-  w(  �  q(  q(   lt 	��1  w(  �  q(  q(   ��  	eF  ~   �  ~(  ~(  �   �K  	�9  �  �  ~(   �(  	
!  ~(    ~(  �  q(   1  	�A  �(  )  �(  ~(  �   �5  	�'  �(  M  �(  ~(  �   �3  	�A  �(  q  �(  �  4   +  	:  4  �  �(   ?  �C  	 �P  ?  �  q(   �B  	$6  w(  �  �(  �(   eof 	(�:  ?  ?  	,N0  ?  �(    _� 
�7   
5�(  
6�)  
7�)  �?  
�%   K  \�  �$   �e  _�  �4  c�)  �J  d�)  ��  qb  h  *   ��  sx  �  *  *   W  y�  *  ~       �J  p  �B  �     %  �   �B  �  $*  �  *    �e  y.  [V    �  �G  !�   <  x  �4  {:  �J  |F  �J  &  `S  �8(  ~J  �  �J  �  �%  ��  �K  ��   I  ��  :!  ��)   %H  �M  h   �3  2  �G  7�  t3  BN*   �'  ��O  <*  !V  ��N  w(  �  �  Y*   !3  �o+  w(      Y*   "�P  ��O  (  .  6*   "�M  ��P  A  G  6*   "�,  �-  Z  e  6*  �   !�+  ��R  �  |  �  6*   !3  �   �  �  �  6*  *  *   �/  !�B  6*  �  �  �  *   "�O  �|6  �  �  6*  *   #(  ��6  �  
  6*  *   $�   �-  �  "  (  6*   %�1  o�*  �  <  6*  *  �    $�A  $n%  �  e  k  **   $�A  (�I  �  �  �  0*  �   $"A  ,�%  6*  �  �  **   $�1  2E)  8  �  �  **   $�/  6;&  8  �  �  **   #�>  :�>  �    0*   $S  A:2  �    *  **  �  �   #�#  K�(  >  S  **  �  �  �   $9  S>$  �  k  {  **  �  �   $-U  [�7  w(  �  �  **  �   &�5  d�-  �  �  �  �   &	1  m�P  �  �  �  �   &�3  v\-  �  �  �  >    &nU  ��-  	  �  8  8   &nU  �nG  >	  �  D  D   &nU  ��   ^	  �  �  �   &nU  �IP  ~	  �  �  �   �J  �rR  ~   �	  �  �   #�=  ��H  �	  �	  0*  �  �  �   #V  �)  �	  �	  0*   '�'  �D*  <*  (�0  �
  
  0*   )�0  �
  "
  0*  *   �0  �2
  =
  0*  B*   �0  �M
  b
  0*  B*  �  �   �0  �r
  �
  0*  B*  �  �  *   �0  ��
  �
  0*  �  �  *   �0  ��
  �
  0*  �  *   �0  ��
  �
  0*  �  >   *   (�0  "    0*  ~    *�  *,Q  H*  +  6  0*  B*   *�  2�G  H*  O  Z  0*  �   *�  =�%  H*  s  ~  0*  >    *S� f�&  8  �  �  0*   *S� q�>  D  �  �  **   +end y<  8  �  �  0*   +end �6;  D  �  �  **   *I ��$  \      0*   *I ��7  P  2  8  **   *��  �lC  \  Q  W  0*   *��  �CM  P  p  v  **   *r ��R  �  �  �  **   *�K  �r5  �  �  �  **   *�3  �j=  �  �  �  **   ,�� �  �  �  0*  �  >    ,�� ��F      0*  �   *I  v  �  1  7  **   ,�E  �|U  L  W  0*  �   ,�1  -�  l  r  0*   *�� 5�?  w(  �  �  **   *�:  D�6  ,  �  �  **  �   *�:  UW     �  �  0*  �   +at k
/  ,  �  �  **  �   +at ��7         0*  �   *�F  ��/  H*  8  C  0*  B*   *�F  �k:  H*  \  g  0*  �   *�F  ��H  H*  �  �  0*  >    *@  DA:  H*  �  �  0*  B*   *@  U�1  H*  �  �  0*  B*  �  �   *@  )�D  H*  �    0*  �  �   *@  ��*  H*    *  0*  �   *@  �6  H*  C  S  0*  �  >    ,�G  -aN  h  s  0*  >    -�3  �b*  H*  �  �  0*  B*   *�3  ^ 2  H*  �  �  0*  B*  �  �   *�3  �=  H*  �  �  0*  �  �   *�3  z�T  H*      0*  �   *�3  � @  H*  *  :  0*  �  >    ,� ��E  O  d  0*  8  �  >    *� �\+  H*  }  �  0*  �  B*   *� �u>  H*  �  �  0*  �  B*  �  �   *� g|=  H*  �  �  0*  �  �  �   *� "�@  H*      0*  �  �   *� 9k<  H*  0  E  0*  �  �  >    *� K�'  8  ^  n  0*  8  >    *bL  d�R  H*  �  �  0*  �  �   *bL  t�2  8  �  �  0*  8   *bL  �L&  8  �  �  0*  8  8   *�%  �9F  H*  �    0*  �  �  B*   *�%  �|<  H*  +  J  0*  �  �  B*  �  �   *�%  ��T  H*  c  }  0*  �  �  �  �   *�%  ��A  H*  �  �  0*  �  �  �   *�%  b>  H*  �  �  0*  �  �  �  >    *�%  3%  H*  �    0*  8  8  B*   *�%  'V7  H*  %  ?  0*  8  8  �  �   *�%  <�+  H*  X  m  0*  8  8  �   *�%  Q'S  H*  �  �  0*  8  8  �  >    *�%  vj.  H*  �  �  0*  8  8  �  �   *�%  ��9  H*  �    0*  8  8  �  �   *�%  �C  H*    9  0*  8  8  8  8   *�%  �>/  H*  R  l  0*  8  8  D  D   $�?  ��&  H*  �  �  0*  �  �  �  >    $�1  �O  H*  �  �  0*  �  �  �  �   ,)  �z-  �  �  �  >   *   .+E  �3J  �    �  >   *   *�5  ��)  �  0  E  **  �  �  �   ,n	 @D  Z  e  0*  H*   *W�  �6  �  ~  �  **   *�A  %�A  �  �  �  **   *��  ,Z5    �  �  **   *�(  �;  �  �  �  **  �  �  �   *�(  I�%  �  	    **  B*  �   *�(  X�5  �  2  B  **  �  �   *�(  �^   �  [  k  **  >   �   *�(  v�S  �  �  �  **  B*  �   *�(  	K  �  �  �  **  �  �  �   *�(  �o?  �  �  �  **  �  �   *�(  J5  �      **  >   �   *NW  ��Q  �  -  =  **  B*  �   *NW  /�I  �  V  k  **  �  �  �   *NW  ��,  �  �  �  **  �  �   *NW  ��;  �  �  �  **  >   �   *�S  ��I  �  �  �  **  B*  �   *�S  >T?  �  �    **  �  �  �   *�S  05  �  -  =  **  �  �   *�S  $S:  �  V  f  **  >   �   *�>  2hL  �    �  **  B*  �   *�>  SUB  �  �  �  **  �  �  �   *�>  Q�2  �  �  �  **  �  �   *�>  _�K  �  �    **  >   �   *�4  qT  �  (  8  **  B*  �   *�4  j�K  �  Q  f  **  �  �  �   *�4  ��5  �    �  **  �  �   *�4  N.  �  �  �  **  >   �   *U+  �)  �  �  �  **  �  �   *��  �!1  ~   �    **  B*   *��  ��T  ~     3  **  �  �  B*   *��  ��O  ~   L  k  **  �  �  B*  �  �   *��  �;.  ~   �  �  **  �   *��  ��B  ~   �  �  **  �  �  �   *��  ��,  ~   �  �  **  �  �  �  �   �  /!T  >   0�E  (  0�F     1�&  1�7  �  �o  >�   �| C~   2Q  bE   ,  2�F cE  2�R  dE  23  eE  2�  fE  2�K  gE  2�@  hE   3all iE  ?4�� ��  :!  ��)   NF  ��*  �E  ��  p0  ��*  �%  ��*  5S  ��*  5�R  ��*  53  ��*  5�$  ��*  5�K  ��*  5�@  ��*  5�@  ��*  #�4  �Z  \  b  _*   #�=  y)  v  |  _*   6�� �  �  _*  �*  �   6�� �  �  _*  �  �   6�� �  �  _*  �   6N  �  �  _*  ~    6��     _*  �*   #�  �U  !  ,  _*  �*   $�&  �.  w(  D  J  _*   #�F  &�;  ^  n  _*  �*  ,   #�9  )�Q  �  �  _*  �*  �*   #WR  ,`2  �  �  _*  �*  �*   #�S  /=  �  �  _*  �*  �*   7e  7,  �  _*  �*  �    �$  _*   5OD  _*  5gP  _*  5�F  $e*  1< 8id ��  �U  ��   5�I  ��)  #�  �<?  k  v  �*  �*   9id ��  �  �*  �*   :id ��  �  �*   ;4H  ��(  �  �  �*    �o  u�  �  u*   �o  ~�  �  u*  {*   )�o  �    u*  �   �o  �  3  u*  {*  �  ,   �o  �C  X  u*  {*  {*  ,   5  �h  s  u*  ~    -�  ��*  {*  �  �  u*  {*   -H�  ��N  �   �  �  �*   -U  �9  w(  �  �  �*  {*   -2  �t*  w(  �  �  �*  {*   <jP  �D        {*   =RD  �Q  {*  >�o  76   A   u*  _*   ?�K  :�N  ?�A  =�5  �K  @I  ,  s   ,   #�,  CH<  �   �   u*  {*  {*  ,   1  ,  �      � >�  @W  3K!  A�4  A�$  Aq-  Ac=  Ao'  A�5   A�%  � A�8  �AX)  �A�%  �A�  �AaO  �AY=  � AP  �� A�C  ��AwS  �A�O  � A�?  �A�5  �� @
$ g�!  A)W  A�   A�U  A�A  A�8  A�P   AEH  �� @�4  ��!  AO   A�7  A(  A�Q  AG  �� Bb4 �#  C�3 ��!  A�3  Ax0 AC5  Df3 &�, �!  �!  �,   -�= 1�,    "  "  �,  {*   �P  ��   E�4  2"  "  Fdec 2"  Et-  2"  Fhex 2"  Er'  2"  E< 2"   Foct 2"  @E� 2"  �G[)  2"   G�%  "2"   G�  &2"   GdO  )2"   G\=  ,2"   G�P  /2"    G�C  32"   @EzS  62"  �E�O  92"  JG�?  <2"  H�  J�!  E�7  NH#  -#  E(  QH#  E�Q  VH#  EO  YH#   H�9  iK!  Fin w�#  w#  Fout z�#  I8- �'3 �#  �,  �!    
<�*  
=�*  
>�*  
@~+  
A�+  
B�+  
C�+  
D�+  
E�+  
F,  
G.,  
HC,  ד  �L$  ��  �  � ��  �4  ��)  /{�  �   J�*  O�   �   �     K$   �C(  �  $
,�  
-  K  :&  �e  =�  � ?�  "  @�  �4  A�)  �J  B�)  �A  O�$  �$  �)   �A  Q�$  �$  �)  *   �A  V%  %  �)  ~    -�
 Y51  �$  /%  :%  *  �$   -�
 ]�R  �$  R%  ]%  *  �$   -� c?  �$  u%  �%  �)  �$  �   D_ m.   �%  �%  �)  �$  �$   -�3  q89  �$  �%  �%  *   D.E  ��3  �%  �%  �)  �$  �)   D�(  ��(  �%  
&  �)  �$   L_Tp >    �$  MZD  �8(  NF�  ��   H��  �!$  H�4  �7$  H� �,$  (��  �l&  r&  g,   O��  ��&  �&  g,  m,   **  ��}  A&  �&  �&  x,   *Ư  �?s  N&  �&  �&  x,   *�F  �Ϭ  ~,  �&  �&  g,   *�F  ��  &  '  '  g,  ~    *a�  �
�  ~,  ('  .'  g,   *a�   ��  &  G'  R'  g,  ~    *�:  ,�  A&  k'  v'  x,  4&   *�F  		n  ~,  �'  �'  g,  4&   *(*  ��  &  �'  �'  x,  4&   * I  h�  ~,  �'  �'  g,  4&   *�O  7k  &  �'  (  x,  4&   *WC  ]�  m,  (  %(  x,   /{�  �  /�  �   18E  &   �� �� �� K2*  7k(  P8!   Q4  Qd  �  d  4  Q�  �  8�)  �{  �   ]�  �  \�   �  �D  !�  �3  "�  U>  #�  &�  $�  �  %�  �*  &�   ڡ  '>   $�U  (>   %TL  )>   &�I  *>   'Q  +>   (�C  ,>   )�J  ->   *1  .�  ,o(  />   0�U  0>   1PL  1>   2�I  2>   3Q  3>   4�C  4>   5�J  5>   6 R)%  K�  �)  ~   �   SGT  P�)  �(  �   ~   Q>   Q�  �$  Q&  &    Q�    �    �  �  Q�  Q  Q�  T7   Y*  U �  �  j*  p*  �     Q�   �   1  Q�   �   �*  �   �  T�*  �*  U T�*  �*  U �*  �*  Q�   �   �l  %   j�  #%   Vtm ,,~+  ,g  .~    �  /~   �  0~   ��  1~   ��  2~   ��  3~   ��  4~   �  5~   d�  6~    ��  7%   $~�  8�  ( S\�  >�*  Rѯ  HJ(  �+  �*  �*   R��  M�*  �+  �+   �*  R�  C�*  �+  �+   �*  R#�  a�  �+  �+   �+  �*  R�� f�  ,  ,   ,  �*  R��  W�+  .,  ,   R[v  \�+  C,  ,   R��  R,   g,  �  ,   �  �+   &  Qs,  �  =(  Q&  WL$  �,  X__a O�   X__b O�    �!  Y�!  �B   ��,  �,  Zh  �,  � [�\�s  [� �,  Y�!  �9   ��,  I-  Zh  �,  �]ȱ  1I-  �^�&   _'U  3   � [�\�s  \��#    {*  `U  =Z-   �   `�   >Z-  `B  ?Z-  `�  E�-   �   `B   F�-  `C  G�-  `e  H�-  `8  I�-  `�  J�-  `

  X�-   �   `�  Y�-  `�
  Z�-  a�   `�-  �   `�  f
.   �   `�  g
.  `�  h
.  `�  n3.   �   `�	  o3.  `�  p3.  `H  v\.   �   ``  w\.  `w  x\.  `   y\.  `~  �.   �   `   ��.  `�  ��.  `  ��.  `�   ��.  `�  ��.  `�	  ��.  `�  ��.   �   `  ��.  `  ��.  `�  ��.  `�  �/     `�  �/  `�  �/  `�  �/  `m  �T/     `	  �T/  `2	  �T/  `�  �T/  `9  �T/  `[  ��/     `J  ��/  `�  ��/  `7  ��/  `�  ��/   "  `I	  ��/  `$	  ��/  `�   ��/   -  `N  ��/  `p  �0   8  `�  �0  `:  �0  `�  �0  `d   �0  `�  �Q0   C  `  �Q0  `�  �Q0  `�	  �z0   N  `�  �z0  `  ؗ0   Y  `�  ٗ0  `�  ڗ0  `�  ۗ0  `+  ��0   d  `�  ��0  `�   ��0  `  ��0   o  `�
  ��0  `�  ��0  `  �1   z  `   �1  `F  �1  `�  �G1   �  `�  �G1  `�  �G1  `D  Op1   �  `�  Pp1  `1  Qp1  `�  W�1   �  `^  X�1  `�  3�1   �  `�  4�1  `�   8�1   �  `�  9�1  `l	  =�1  �  `N  >�1  `^  ?�1  `L  @�1  `a  D%2  �  `B  E%2  `�	  F%2  `  G%2  `  H%2  `y  I%2  `�   r2   �  `�  !r2   R    * K� �� �V  �F     �� �  (  _� �>   �  �  P   �  �  o  �	  pW   w   �  qW  !�   int   "�   �    #�   #  s  NE   �  VE   Fd ~   Z�  l   .  <~   `  D�   �  W~   �  _�   �  e�   t   m�   a  u�     ~�   �  ��   3  ��   �  ��   H  ��   y  ��     ��   s  ��   T   ȉ   �  Љ   F  ׉   �  ��   �  �     �   V  �   %   �  \	  2�   o  7�   �  <�   �  C�   �  �   E   	\  �   gX  �   � �   <�  �   B� #�   � $�   E� %�   � &�   Q� '�   X\  	&�  X\  X	,�  	$Z  	.�    	\ 	/E   	� 	1  	Z  	23   	K]  	3E   	�_  	43   	\W  	53   	�Z  	63   	-_  	8�   	VY  	9�  $	`  	:  (	�Y  	;  ,	7_  	<.  0	BY  	=X  4	b\  	>.  8	\  	?.  <	7Y  	@.  @	 Z  	Ai  D	SX  	Bi  H	n4 	Dl   L	`  	F�  P	*5 	G�  T 
(  �  �   3   �   �  �  
(  �  �  3   �   �  �  
�     �    �    �  
    �   
  
�   .  �     
�  M  M  M  �   S  %   4  i  �   ^  �^  
!  std  �  b�  co  e�  f�  g  h)  i?  jT  kj  l�  m�  q�  r�  t	  u)  vO  xe  y{  |�  ~�  ��  ��  ��  ��  �  �)  �4  �I  @w  %  0�:  Z�   _� �>   5�  6�  7  �?  �,   W  3  �4  �$  q-  c=  o'  �5   �%  � �8  �X)  ��%  ��  �aO  �Y=  � P  �� �C  ��wS  ��O  � �?  ��5  �� 
$ gU  )W  �   �U  �A  �8  �P   EH  �� �4  ��  O   �7  (  �Q  G  �� ��  ��  �R   �-  �1  lO  �� b4 �  �9  i  �N  ��  �P  ��  �4  �  �  dec �  t-  �  hex �  r'  �  < �   oct �  @� �  �[)  �   �%  "�   �  &�   dO  )�   \=  ,�   �P  /�    �C  3�   @zS  6�  ��O  9�  J�?  <�  �  JU  �7  N�  �  (  Q�  �Q  V�  O  Y�   app l9  �  @� t9  in w9  out z9  �P  }9   cur ��  �   �  5�
  	 8;   	��  ;�  � >�  �  A  G   @�  Ad�  A  �  �  A  M  �  �    &�  Dx�  A  	  	  A  ;  �   &�  G( A  5	  E	  A  �   �   <_  JG�  A  ]	  c	  A   �  M��  �  {	  �	  M   fd P� �   �	  �	  A   QY  S� ;  �	  �	  A   � U�	  �	  A  �    �W  X" �
  �	  �	  A  M  �
   f [� �
  
  1
  A  M  �
  M  �
   �W  _: �
  I
  Y
  A  �  �
   09  b��  W  q
  �
  A  W  �   � e  �   �
  �
  A   ��  h��  �
  �
  A    �^  -�  � *d  �  �>  b�  �0 �  R1 �1  �1 �2 �3  F2 �*  / v/  �4    �
   �� ��  !�+ �6  !}�  �1  ?!�. �1  !�3 6  !�. 6  !J- 6  !_5 1  !�4 1   !r6 1   !f1 1   !0 1   !/, 6   !�1 6   !Y2 6   !V, *   !5 6   !x, '6   !�+ (6  !�2 )6   !�4 +6  !�3 ,6   !�0 -/   "min ��� �   "max ��� �   #T4 	�� �   #/5 � �   #�2 �� �   #�1 �� �   #]2 !'� �   #�4 %J� �    �
   $Z  
1�  �   �  %aY  
��     �   &\  
C�   )  �   &xZ  
M�   ?  �   %`  
��   T  �   &�^  
r�   j  �   &_X  
��   �  �  �   o  &�_  
��  �  �  �   �   %�\  
��  �  M  M   &4Z  
�3   �  �  3   3   �   %7`  
��  	  M  M  �   &>]  
	�   )  �  ,   �    &�Z  
�   D  �  D   J  o  &�Y  
 ,   e  �   &�Y  
��   {  �   '\  
��   %�_  0�  �  �   $�]  
W�  M   %D[  
T�   �  M   %�[  
a�   �  M  M   $�\  
)�  �   (Y@ 
�  �  �   %�[  
   )  �  �  �   3    )�]  
i�  %D]  
w�  I  �   &}W  
��   d  �   �   ��  !�   *pO qO !o  +$   ��  �  $,b  -�   �� �� �� +2*  7�  ,8P   �  �  8�  	�{  �   	]�  �  	\�   �  	�D  !�  	�3  "�  	U>  #�  	&�  $�  	�  %�  	�*  &�   	ڡ  '%   $	�U  (%   %	TL  )%   &	�I  *%   '	Q  +%   (	�C  ,%   )	�J  -%   *	1  .�  ,	o(  /%   0	�U  0%   1	PL  1%   2	�I  2%   3	Q  3%   4	�C  4%   5	�J  5%   6 %)%  K�    �   M   )GT  P$  �    �   �  �
  �  �
  �
  c� l   �l  ,   � 42  	y� 4>   	>� 53  	� 6S  	�� 7I  	�� 8T  	�� 9_  	� :  	j� ;^   	�� <^  $	�� =^  (	�� >j  ,	�� ?u  0 -<  .q� IM     �   /�� r�
  �   M  �
    ,E  0  Z  1�% I�  2 3c	  �j  t  4h  t   M  5o  5_  6�
  L�  �  4h  �   A  7   S   �  8� r�   �� 9__s rM  �� 9__n r�
  �� :`E ;�s t�
  �� :�E ;�&  x�  #� <A�     3�  � )  8  4h  �  G   =  �� p   �S  d  >)  � >2  � ?�  ��f   �}  �  @h  �  � A
� �;  �B�  �:�E ;�&  �A  A� C�@   ;�*  Ɖ   x� D�  �	   �E�  �� <�?      ?	  ���   �	  �  @h  �  � A� ։   �A^F  ֲ  �F�E �  ;�&  �A  �� G�� �M  HC  ��E �v  EM  �� I�E  F�E �  ;��  ��  %� <\   <<�   <t�  <}�   ?�  �Q   ��  I  @h  �  � AF�  �M  �A^F  �  �B�   �:F ;�&  �A  9� G�� �M  HC  �@F �>  >M  �I@F  <��    =Z  ��  �   �d  m  >j  �  ?�	  ��,   ��  �  @h  �  � < �  <�  <�   J�	      ��  �  @h  �  �  JE	  0n   ��  O  @h  �  � :XF K�&  	A  z� LZ  9   
.  Ej  ��  :�F K�*  �   �� <v�     3�	  � _  r  4h  �  4#  1   =O  !� �   ��  �  >_  � M��  N� �   J1
   �Q   ��    @h  �  � O__s  �  �O__n  �
  �:�F K�&  "�
  )� <�m  <��    J�	  *$   �/  {  @h  �  � O__s *M  �O__n *�
  �<&m  M4�  NR�NQ�  J�	  .@h   ��  9  @h  �  � P�e  .M  �P7i .�
  �P�e  /M  �P<i /�
  �:�F K�&  1�
  G� <[m  Qk�    NR�NQ� <�m  R��  NR�NQv    JY
  ?�E   �S  �  @h  �  � PQ  ?W  �P@  ?�  �<�m  <�  <��  <��   =�        ��  �  E�  �� S?   J�
  PP   ��  E  @h  �  � C?   T� qi  ��K�*  r1  �� <m  <,5  <Bm  <Q    UD  OQ   �   U�  PQ  U1  QQ  U�  Wz   �   U^  Xz  UU  =�   �   U�   >�  UB  ?�  U�  E�   �   UB   F�  UC  G�  Ue  H�  U8  I�  U�  J�  U

  X   �   U�  Y  U�
  Z  V�   `6    U�  fG     U�  gG  U�  hG  U�  np     U�	  op  U�  pp  UH  v�   #  U`  w�  Uw  x�  U   y�  U~  �   .  U   ��  U�  ��  U  ��  U�   ��  U�  ��  U�	  ��  U�  �'   9  U  �'  U  �'  U�  �'  U�  �\   D  U�  �\  U�  �\  U�  �\  Um  ��   O  U	  ��  U2	  ��  U�  ��  U9  ��  U[  ��   Z  UJ  ��  U�  ��  U7  ��  U�  �   e  UI	  �  U$	  �  U�   �0   p  UN  �0  Up  �M   {  U�  �M  U:  �M  U�  �M  Ud   �M  U�  Ɏ   �  U  ʎ  U�  ˎ  U�	  ѷ   �  U�  ҷ  U  ��   �  U�  ��  U�  ��  U�  ��  U+  �	   �  U�  �	  U�   �	  U  �2   �  U�
  �2  U�  �2  U  �[   �  U   �[  UF  �[  U�  �   �  U�  �  U�  ��  U�  3�   �  U�  4�  U�   8�   �  U�  9�  Ul	  =�  �  UN  >�  U^  ?�  UL  @�  Ua  D    UB  E  U�	  F  U  G  U  H  Uy  I  U�   i     U�  !i  W|�  �   %�9  .(  �  �   �  3    &�� 
j�  �  �   M   X>  Y  �  �    Y  �  �    &g\  
a�   �  �   %2_  )(    �   �   3    %s� 3  5  �     �    %� F�   O  �   O   i   g)   �. �� m� �V  hG     y� (  _� �7   �  �  8k  �{  k   ]�  k  \�   k  �D  !k  �3  "k  U>  #k  &�  $k  �  %k  �*  &k   ڡ  'q  $�U  (q  %TL  )q  &�I  *q  'Q  +q  (�C  ,q  )�J  -q  *1  .k  ,o(  /q  0�U  0q  1PL  1q  2�I  2q  3Q  3q  4�C  4q  5�J  5q  6 q  �  std  �  5>   6�  7�  @u  	%  0�=  �n  �b  �q  Fe  �  
�3  �=  �  �!  �!   �  eq �<-  �!    �!  �!   lt ��1  �!  !  �!  �!   ��  eF  �  E  �!  �!  n   �K  �9  n  _  �!   �(  
!  �!  �  �!  n  �!   1  �A  �!  �  �!  �!  n   �5  �'  �!  �  �!  �!  n   �3  �A  �!  �  �!  n  �   +  :  �  	  �!   �  �C   �P  �  (  �!   �B  $6  �!  G  �!  �!   eof (�:  �  ?  ,N0  �  �!    _� �7   �?  �%   K  \  �   �e  _n  �4  c�!  �J  d�!  ��  q�  �  �!   ��  s�  �  �!  �!   W  y�  �!  �    �  �J  	pz  �B  	R  �   %  	k   �B  	A  �!  k  �!    �e  	y�  [V  	k  R  �G  	!   <  	x�  �4  	{�  �J  	|�  �J  	6  `S  	�U!  ~J  	�z  �J  	�  �%  	�  �K  	�R   I  	�R  :!  	��!   %H  	��  �   �3  
2k  �G  
7�  t3  
B"  �'  	��O  "  V  	��N  �!  [  a  "   3  	�o+  �!  x  ~  "   �P  	��O  �  �  �!   �M  	��P  �  �  �!   �,  	�-  �  �  �!  R   �+  	��R  k  �  �  �!   3  	�   k      �!  �!  �!   �/  
!�B  �!  6  R  R  �!   �O  	�|6  I  T  �!  �!    (  
��6  h  s  �!  �!   !�   	�-  k  �  �  �!   "�1  
o�*  k  �  �!  �!  R    !�A  	$n%  k  �  �  �!   !�A  	(�I  k  �  �  �!  k   !"A  	,�%  �!      �!   !�1  	2E)  �  -  3  �!   !�/  	6;&  �  K  Q  �!    �>  	:�>  e  k  �!   !S  	A:2  R  �  �  �!  R  �    �#  	K�(  �  �  �!  R  R  �   !9  	S>$  R  �  �  �!  R  R   !-U  	[�7  �!  �    �!  �   #�5  	d�-  '  k  �  R   #	1  	m�P  G  k  �  R   #�3  	v\-  g  k  R  q   #nU  	��-  �  k  �  �   #nU  	�nG  �  k  �  �   #nU  	��   �  k  k  k   #nU  	�IP  �  k  �  �   �J  	�rR  �  	  R  R    �=  
��H  	  /	  �!  R  R  R    V  
�)  C	  I	  �!   $�'  	�D*  "  %�0  	�j	  p	  �!   &�0  
��	  �	  �!  �!   �0  
��	  �	  �!  "   �0  
��	  �	  �!  "  R  R   �0  
��	  �	  �!  "  R  R  �!   �0  
�
  
  �!  �  R  �!   �0  
�*
  :
  �!  �  �!   �0  
�J
  _
  �!  R  q  �!   %�0  	"p
  {
  �!  �   '�  	*,Q  "  �
  �
  �!  "   '�  	2�G  "  �
  �
  �!  �   '�  	=�%  "  �
  �
  �!  q   'S� 	f�&  �       �!   'S� 	q�>  �    %  �!   (end 	y<  �  >  D  �!   (end 	�6;  �  ]  c  �!   'I 	��$  �  |  �  �!   'I 	��7  �  �  �  �!   '��  	�lC  �  �  �  �!   '��  	�CM  �  �  �  �!   'r 	��R  R  �  �  �!   '�K  	�r5  R      �!   '�3  	�j=  R  6  <  �!   )�� 
�  Q  a  �!  R  q   )�� 	��F  v  �  �!  R   'I  	v  R  �  �  �!   )�E  
�|U  �  �  �!  R   )�1  	-�  �  �  �!   '�� 	5�?  �!  �  �  �!   '�:  	D�6  �      �!  R   '�:  	UW  �  7  B  �!  R   (at 	k
/  �  Z  e  �!  R   (at 	��7  �  }  �  �!  R   '�F  	��/  "  �  �  �!  "   '�F  	�k:  "  �  �  �!  �   '�F  	��H  "  �  �  �!  q   '@  
DA:  "      �!  "   '@  
U�1  "  1  F  �!  "  R  R   '@  
)�D  "  _  o  �!  �  R   '@  	��*  "  �  �  �!  �   '@  
�6  "  �  �  �!  R  q   )�G  	-aN  �  �  �!  q   *�3  
�b*  "  �  �  �!  "   '�3  	^ 2  "    -  �!  "  R  R   '�3  
�=  "  F  V  �!  �  R   '�3  	z�T  "  o  z  �!  �   '�3  	� @  "  �  �  �!  R  q   )� 	��E  �  �  �!  �  R  q   '� 	�\+  "  �  �  �!  R  "   '� 	�u>  "    )  �!  R  "  R  R   '� 
g|=  "  B  W  �!  R  �  R   '� 	"�@  "  p  �  �!  R  �   '� 	9k<  "  �  �  �!  R  R  q   '� 	K�'  �  �  �  �!  �  q   'bL  	d�R  "  �     �!  R  R   'bL  	t�2  �    $  �!  �   'bL  
�L&  �  =  M  �!  �  �   '�%  	�9F  "  f  {  �!  R  R  "   '�%  	�|<  "  �  �  �!  R  R  "  R  R   '�%  
��T  "  �  �  �!  R  R  �  R   '�%  	��A  "  �    �!  R  R  �   '�%  	b>  "  -  G  �!  R  R  R  q   '�%  	3%  "  `  u  �!  �  �  "   '�%  	'V7  "  �  �  �!  �  �  �  R   '�%  	<�+  "  �  �  �!  �  �  �   '�%  	Q'S  "  �  	  �!  �  �  R  q   '�%  	vj.  "  "  <  �!  �  �  k  k   '�%  	��9  "  U  o  �!  �  �  �  �   '�%  	�C  "  �  �  �!  �  �  �  �   '�%  	�>/  "  �  �  �!  �  �  �  �   !�?  
��&  "  �    �!  R  R  R  q   !�1  
�O  "    9  �!  R  R  �  R   ,)  	�z-  k  ]  R  q  �!   ++E  
�3J  k  �  R  q  �!   '�5  
��)  R  �  �  �!  k  R  R   )n	 
@D  �  �  �!  "   'W�  	�6  �  �  �  �!   '�A  	%�A  �      �!   '��  	,Z5  }  %  +  �!   '�(  
�;  R  D  Y  �!  �  R  R   '�(  	I�%  R  r  �  �!  "  R   '�(  	X�5  R  �  �  �!  �  R   '�(  
�^   R  �  �  �!  q  R   '�(  	v�S  R  �  �  �!  "  R   '�(  
	K  R    +  �!  �  R  R   '�(  	�o?  R  D  T  �!  �  R   '�(  
J5  R  m  }  �!  q  R   'NW  	��Q  R  �  �  �!  "  R   'NW  
/�I  R  �  �  �!  �  R  R   'NW  	��,  R  �  �  �!  �  R   'NW  	��;  R    &  �!  q  R   '�S  	��I  R  ?  O  �!  "  R   '�S  
>T?  R  h  }  �!  �  R  R   '�S  	05  R  �  �  �!  �  R   '�S  	$S:  R  �  �  �!  q  R   '�>  	2hL  R  �  �  �!  "  R   '�>  
SUB  R    &  �!  �  R  R   '�>  	Q�2  R  ?  O  �!  �  R   '�>  
_�K  R  h  x  �!  q  R   '�4  	qT  R  �  �  �!  "  R   '�4  
j�K  R  �  �  �!  �  R  R   '�4  	��5  R  �  �  �!  �  R   '�4  
N.  R    !  �!  q  R   'U+  	�)  	  :  J  �!  R  R   '��  	�!1  �  c  n  �!  "   '��  
��T  �  �  �  �!  R  R  "   '��  
��O  �  �  �  �!  R  R  "  R  R   '��  
�;.  �  �  �  �!  �   '��  
��B  �    &  �!  R  R  �   '��  
��,  �  ?  Y  �!  R  R  �  R     ,!T  q  -�E  �  -�F  �   .�&  .�7  	  � >	  </"  =$"  >:"  @�"  A�"  B�"  C
#  D%#  EE#  Fe#  Gz#  H�#  ۝  �  /@�  ��   ד  �9  ��  �y  � �k  �4  ��!  ,{�  k   0l�  �  1�  (Uo  �  9  b  |  �#  �  �  �  �#   ,!T  q   9  �   2)%  Kk  �  �  �   3int �  q  4GT  P�  >   �  �  �  �  o  �	  �  qW  !�    "  �  #  .  <�  `  D�  �  W�  �  _  �  e�  t   m�  a  u�    ~�  �  ��  3  ��  �  ��  H  ��  y  ��    ��  s  ��  T   ȫ  �  Ы  F  ׫  �  �  �  �    �  V  �  �  s  N�  �  V�  \	  2�  o  7�  �  <�  �  C�  �  �  l  56pO qO !m  7$   E`!  	�  $,n  -y  K  :1  �e  =n  � ?k  "  @�  �4  A�!  �J  B�!  �A  O�  �  �!   �A  Q    �!  �!   �A  V)  4  �!  �   *�
 Y51  �  L  W  �!  �   *�
 ]�R  �  o  z  �!  �   *� c?  �  �  �  �!  �  f   8_ m.   �  �  �!  �  �   *�3  q89  �  �  �  �!   8.E  ��3  �    �!  �  �!   8�(  ��(    '  �!  �   9_Tp q   �  :ZD  �U!  ;F�  �k   <��  �  <�4  �$  <� �  %��  ��  �  �#   =��  ��  �  �#  �#   '*  ��}  ^  �  �  �#   'Ư  �?s  k  �  �  �#   '�F  �Ϭ  �#        �#   '�F  ��  6  !   ,   �#  �   'a�  �
�  �#  E   K   �#   'a�   ��  6  d   o   �#  �   '�:  ,�  ^  �   �   �#  Q   '�F  		n  �#  �   �   �#  Q   '(*  ��  6  �   �   �#  Q   ' I  h�  �#  �   �   �#  Q   '�O  7k  6  !  #!  �#  Q   'WC  ]�  �#  <!  B!  �#   ,{�  k  ,�  	   .8E  6   �� �� �� 72*  7�!  >8�   ?�  ?�  �  �  �  ?	  ?q  ?�  �  ?1  1  �  ?    �   �    �  	    ?  ?�  ?	  @7   "  A Y  �l  %   j�  #%   Btm ,,�"  ,g  .�   �  /�  �  0�  ��  1�  ��  2�  ��  3�  ��  4�  �  5�  d�  6�   ��  7%   $~�  8�  ( 4\�  >/"  2ѯ  Hg!  �"  $"  $"   2��  M$"  #  #   :"  2�  C$"  #  #   $"  2#�  ak  :#  :#   @#  :"  2�� fk  Z#  Z#   `#  $"  2��  W#  z#  Z#   2[v  \#  �#  Z#   2��  R,   �#  k  ,   �  :#   6  ?�#  k  Z!  ?6  �  ?�  CB  `   ��#  +$  Dh  +$  �E�  �E�  �E�  �F�  (0$  �Gr �#  �#  HU  =A$      H�   >A$  HB  ?A$  H�  Ej$   +  HB   Fj$  HC  Gj$  He  Hj$  H8  Ij$  H�  Jj$  H

  X�$   6  H�  Y�$  H�
  Z�$  I�   `�$  A  H�  f�$   L  H�  g�$  H�  h�$  H�  n%   W  H�	  o%  H�  p%  HH  vC%   b  H`  wC%  Hw  xC%  H   yC%  H~  x%   m  H   �x%  H�  �x%  H  �x%  H�   �x%  H�  �x%  H�	  �x%  H�  ��%   x  H  ��%  H  ��%  H�  ��%  H�  �&   �  H�  �&  H�  �&  H�  �&  Hm  �;&   �  H	  �;&  H2	  �;&  H�  �;&  H9  �;&  H[  �|&   �  HJ  �|&  H�  �|&  H7  �|&  H�  ��&   �  HI	  ��&  H$	  ��&  H�   ��&   �  HN  ��&  Hp  ��&   �  H�  ��&  H:  ��&  H�  ��&  Hd   ��&  H�  �8'   �  H  �8'  H�  �8'  H�	  �a'   �  H�  �a'  H  �~'   �  H�  �~'  H�  �~'  H�  �~'  H+  �'   �  H�  �'  H�   �'  H  ��'   �  H�
  ��'  H�  ��'  H  �(   �  H   �(  HF  �(  H�  �.(     H�  �.(  H�  �.(  HD  OW(     H�  PW(  H1  QW(  H�  W�(   $  H^  X�(  H�  3�(   /  H�  4�(  H�   8�(   :  H�  9�(  Hl	  =�(  E  HN  >�(  H^  ?�(  HL  @�(  Ha  D)  P  HB  E)  H�	  F)  H  G)  H  H)  Hy  I)  H�   Y)   [  H�  !Y)   �6   n3 �� )� �V  HH     9� std  �  %  0@�!  �=  �  �b  �   Fe  ��  �3  �=  z   �!  �!   	J   
eq �<-  �!  �   �!  �!   
lt ��1  �!  �   �!  �!   ��  eF  �  �   �!  �!     �K  �9    �   �!   �(  
!  �!    �!    �!   1  �A  �!  ?  �!  �!     �5  �'  �!  c  �!  �!     �3  �A  �!  �  �!    J    +  :  J   �  �!   	U   �C   �P  U   �  �!   �B  $6  �!  �  �!  �!   eof (�:  U   ?  ,N0  U   �!    _� ��  �?  ��  K  \�  �   �e  _  �4  c�!  �J  d�!  ��  qc  i  �!   ��  sy  �  �!  �!   W  y�  �!  �    	  5"  61#  7K#  �J  p?  �B       %  -!   �B  �    l#  -!  �!   �B    l#  �    �e  y/  [V  0  	  �G  !�   <  x  �4  {;  �J  |G  �J  j  `S  �o  ~J  �?  �J  �D  �%  ��  �K  �   I  �  :!  �\#   %H  �{  �   �3  	20  �G  	7�!  t3  	B�#  �'  ��O  �#  V  ��N  �!     &  �#   3  �o+  �!  =  C  �#   �P  ��O  V  \  ~#   �M  ��P  o  u  ~#   �,  �-  �  �  ~#     �+  ��R  -!  �  �  ~#   3  �   -!  �  �  ~#  �!  �!   �/  	!�B  ~#  �      �!   �O  �|6      ~#  �!   (  	��6  -  8  ~#  �!    �   �-  -!  P  V  ~#   !�1  	o�*  -!  j  ~#  �!       �A  $n%  -!  �  �  r#    �A  (�I  -!  �  �  x#  -!    "A  ,�%  ~#  �  �  r#    �1  2E)  f  �  �  r#    �/  6;&  f      r#   �>  :�>  *  0  x#    S  A:2    H  X  r#    �!   �#  K�(  l  �  r#      �!    9  S>$    �  �  r#        -U  [�7  �!  �  �  r#  �!   "�5  d�-  �  -!  �!     "	1  m�P    -!  �!     "�3  v\-  ,  -!        "nU  ��-  L  -!  f  f   "nU  �nG  l  -!  r  r   "nU  ��   �  -!  -!  -!   "nU  �IP  �  -!  �!  �!   �J  �rR  �  �       �=  	��H  �  �  x#         V  	�)      x#   #�'  �D*  �#  $�0  �/  5  x#   %�0  	�E  P  x#  �!   �0  	�`  k  x#  �#   �0  	�{  �  x#  �#       �0  	��  �  x#  �#      �!   �0  	��  �  x#  �!    �!   �0  	��  �  x#  �!  �!   �0  	�	  $	  x#       �!   $�0  "5	  @	  x#  �   &�  *,Q  �#  Y	  d	  x#  �#   &�  2�G  �#  }	  �	  x#  �!   &�  =�%  �#  �	  �	  x#      &S� f�&  f  �	  �	  x#   &S� q�>  r  �	  �	  r#   'end y<  f  
  	
  x#   'end �6;  r  "
  (
  r#   &I ��$  �  A
  G
  x#   &I ��7  ~  `
  f
  r#   &��  �lC  �  
  �
  x#   &��  �CM  ~  �
  �
  r#   &r ��R    �
  �
  r#   &�K  �r5    �
  �
  r#   &�3  �j=    �
    r#   (�� 	�    &  x#        (�� ��F  ;  F  x#     &I  v    _  e  r#   (�E  	�|U  z  �  x#     (�1  -�  �  �  x#   &�� 5�?  �!  �  �  r#   &�:  D�6  Z  �  �  r#     &�:  UW  N  �    x#     'at k
/  Z    *  r#     'at ��7  N  B  M  x#     &�F  ��/  �#  f  q  x#  �#   &�F  �k:  �#  �  �  x#  �!   &�F  ��H  �#  �  �  x#      &@  	DA:  �#  �  �  x#  �#   &@  	U�1  �#  �    x#  �#       &@  	)�D  �#  $  4  x#  �!     &@  ��*  �#  M  X  x#  �!   &@  	�6  �#  q  �  x#        (�G  -aN  �  �  x#      )�3  	�b*  �#  �  �  x#  �#   &�3  ^ 2  �#  �  �  x#  �#       &�3  	�=  �#      x#  �!     &�3  z�T  �#  4  ?  x#  �!   &�3  � @  �#  X  h  x#        (� ��E  }  �  x#  f        &� �\+  �#  �  �  x#    �#   &� �u>  �#  �  �  x#    �#       &� 	g|=  �#      x#    �!     &� "�@  �#  5  E  x#    �!   &� 9k<  �#  ^  s  x#          &� K�'  f  �  �  x#  f      &bL  d�R  �#  �  �  x#       &bL  t�2  f  �  �  x#  f   &bL  	�L&  f      x#  f  f   &�%  �9F  �#  +  @  x#      �#   &�%  �|<  �#  Y  x  x#      �#       &�%  	��T  �#  �  �  x#      �!     &�%  ��A  �#  �  �  x#      �!   &�%  b>  �#  �    x#            &�%  3%  �#  %  :  x#  f  f  �#   &�%  'V7  �#  S  m  x#  f  f  �!     &�%  <�+  �#  �  �  x#  f  f  �!   &�%  Q'S  �#  �  �  x#  f  f        &�%  vj.  �#  �    x#  f  f  -!  -!   &�%  ��9  �#    4  x#  f  f  �!  �!   &�%  �C  �#  M  g  x#  f  f  f  f   &�%  �>/  �#  �  �  x#  f  f  r  r    �?  	��&  �#  �  �  x#             �1  	�O  �#  �  �  x#      �!     ,)  �z-  -!  "       �!   *+E  	�3J  -!  E       �!   &�5  	��)    ^  s  r#  -!       (n	 	@D  �  �  x#  �#   &W�  �6  �!  �  �  r#   &�A  %�A  �!  �  �  r#   &��  ,Z5  B  �  �  r#   &�(  	�;    	    r#  �!       &�(  I�%    7  G  r#  �#     &�(  X�5    `  p  r#  �!     &�(  	�^     �  �  r#        &�(  v�S    �  �  r#  �#     &�(  		K    �  �  r#  �!       &�(  �o?    	    r#  �!     &�(  	J5    2  B  r#        &NW  ��Q    [  k  r#  �#     &NW  	/�I    �  �  r#  �!       &NW  ��,    �  �  r#  �!     &NW  ��;    �  �  r#        &�S  ��I        r#  �#     &�S  	>T?    -  B  r#  �!       &�S  05    [  k  r#  �!     &�S  $S:    �  �  r#        &�>  2hL    �  �  r#  �#     &�>  	SUB    �  �  r#  �!       &�>  Q�2        r#  �!     &�>  	_�K    -  =  r#        &�4  qT    V  f  r#  �#     &�4  	j�K      �  r#  �!       &�4  ��5    �  �  r#  �!     &�4  	N.    �  �  r#        &U+  �)  �  �    r#       &��  �!1  �  (  3  r#  �#   &��  	��T  �  L  a  r#      �#   &��  	��O  �  z  �  r#      �#       &��  	�;.  �  �  �  r#  �!   &��  	��B  �  �  �  r#      �!   &��  	��,  �      r#      �!     	�  +!T     ,�E  >   ,�F     -�&  -�7  	�  .�{ 
�e  �  �   /�{ s  ~  �#  �#   %�{ T�  �  �#  �#   0�� WN  �  �#  �    .�8 
pe  P  e   K� 
rZ  /�8 �  �  �#  �#   %�8 A    �#  �#   1�� D�  "  -  �#  �   2(� GI� �!  �  I  �#    	N  	Z  � >�  3�� �  �� ?z  �$    .jy 
�e  �  �   /jy �  �  �#  �#   %jy O�  �  �#  �#   0�� R�  �  �#  �    	�  . 
�e  V  �   /     �#  �#   % J.  9  �#  �#   0*� M�  J  �#  �    	�  	�  .�z 
de  �  �   /�z �  �  �#  �#   %�z <�  �  �#  �#   0�� ?`  �  �#  �    .�p 
7e  b  e   K� 
9Z  /�p �    $  $   %�p $    $  �#   1�� '�  4  ?  $  �   2(� *�� �!  �  [  $    	`  .� 
[e  �  �   /� �  �  �#  �#   %� 7�  �  �#  �#   07� :g  �  �#  �    	g  .�� 
Re  <  �   /�� �    �#  $   %�� 2    �#  �#   0�� 5�  0  �#  �    	�  .� 
Je  �  �   /� f  q  $  $   %� -�  �  $  �#   0� 0A  �  $  �    	A  	�   4$   E�  �  $,  -  K  :e  �e  =  � ?-!  "  @�!  �4  A�!  �J  B�!  �A  O,  2  �!   �A  QB  M  �!  �!   �A  V]  h  �!  �   )�
 Y51  �  �  �  �!     )�
 ]�R  �  �  �  �!     )� c?  �  �  �  �!  �  �!   5_ m.   �  �  �!  �  �   )�3  q89  �      �!   5.E  ��3  ,  <  �!  �  �!   5�(  ��(  P  [  �!  �   6_Tp     	�  -ZD  -8E  7U  A\#  �  %$  �   89+  N\#  %$  �    9�  9o  9�  9�  9�  9�  9�	  :int 9(  9#  9�� 9�� 9�� 42*  7   ;80    9�  �  �  qW  !�    "�  .  <%   `  D�  �  W%   �  _0   �  e�  t   m�  a  u�    ~�  �  ��  3  ��  �  ��  H  ��  y  ��    ��  s  ��  T   ��  �  ��  F  ��  �  ��  �  ��    ��  V  ��  <   9�  =s  N   �  V   \	  2�  o  7�  �  <�  �  C�  �  �  <�!  ><�!  	   ?pO qO !�!  @J   @z   9�  <z   <J   @�  @   @�!  <�  @e  <e  <  @�  9  �  81#  �{  -!   ]�  -!  \�   -!  �D  !-!  �3  "-!  U>  #-!  &�  $-!  �  %-!  �*  &-!   ڡ  '   $�U  (   %TL  )   &�I  *   'Q  +   (�C  ,   )�J  -   *1  .-!  ,o(  /   0�U  0   1PL  1   2�I  2   3Q  3   4�C  4   5�J  5   6 A)%  K-!  K#  �  �!   BGT  PV#  <"  �   �  	�  <�  <I  <�  <�  @�  @I  @�  C�  �#  D <  <N  @P  @U  <�  @�  <�  @V  <�  @[  <[  <`  @b  <g  @�  <�  @<  <A  @�  <�  @�  <�  <\#  Et  Y$  FXF  A%$  F\;  A�  GH�T  C\#    I{  g$  q$  Jh  q$   	r#  I�  �$  �$  Jh  q$   E�  �$  GK__p �:!    E�  �$  FXF  N%$  F\;  N�   I�  �$  �$  Jh  �$  L__a ��$   	~#  	�!  <e  In  %  %  Jh  %   	�$  IM  %%  8%  Jh  8%  J#  g#   	�!  I�  K%  ^%  Jh  ^%  J#  g#   	�!  I2  q%  �%  Jh  8%  �%   	�!  Ii  �%  �%  Jh  ^%  L__a s�%   	�!  I�  �%  �%  Jh  q$   I�  �%  �%  Jh  q$   M  �%  &  Jh  &  J#  g#   	l#  I$	  &  '&  Jh  '&  J#  g#   	x#  I�  :&  M&  Jh  M&  J#  g#   	$  I  `&  s&  Jh  s&  J#  g#   	�#  I�  �&  �&  Jh  �&  J#  g#   	�#  I�  �&  �&  Jh  �&  J#  g#   	�#  I9  �&  �&  Jh  �&  J#  g#   	�#  I�  �&  '  Jh  '  J#  g#   	�#  I�  '  1'  Jh  1'  J#  g#   	�#  N?  �   �M'  Z'  Oh  Z'  �  	$  N-  �   �v'  �'  Oh  �'  �  	�#  I   �'  �'  Jh  �'  J#  g#   	$  P�'  E� �P   ��'  �(  Q�'  � R&  �xG '�(  S&  �� T�%  ��G #%(  S�%  �� UY$  �   -Sg$  ��   V�$  ��G #S�$  �� S�$  � W�    S�$  ,� S�$  Y� R�$  ��G ��(  X�$  S�$  l� Y+$  ��G VX@$  S5$  l� Z�G [L$  ��    \�     ]� P,&  � �   ��(  �(  Q:&  � ^��'  _� �   P,&  ��  !   �)  N)  Q:&  � `,&     0D)  S:&  �� \�'   a!�6   PR&  �� 0   �i)  �)  Q`&  � ^?�'  _� �   PR&  y� @!   ��)  �)  Q`&  � `R&  H   5�)  S`&  �� \T�'   aa�6   Px&  �� p   ��)  *  Q�&  � ^�'  _� �   Px&  �� �!   �(*  `*  Q�&  � `x&  �   :V*  S�&  �� \��'   a��6   P�&  � �   �{*  �*  Q�&  � ^��'  _� �   P�&  �� �!   ��*  �*  Q�&  � `�&  �   ?�*  S�&  �� \��'   a��6   P�'  �� �   �+  +  Q�'  � \��'  a�6   I   -+  @+  Jh  @+  J#  g#   	�#  P+  �� P   �`+  \,  Q-+  � R&  �G DV,  S&  � T�%   H #�+  S�%  � UY$     -Sg$  �   V�$  %H #S�$  O� S�$  |� W@    S�$  �� S�$  �� R�$  @0H �J,  X�$  S�$  �� Y+$  @0H VX@$  S5$  �� Z0H [L$  ��    \[     ]6 P�&  �� `   �w,  �,  Q�&  � ^oE+  _� �   P�&  �� p!   ��,  �,  Q�&  � `�&  x   M�,  S�&  � \�E+   a��6   P�&  �� �   � -  -  Q�&  � ^�E+  _� �   P�&  �� �!   �6-  n-  Q�&  � `�&  �   Rd-  S�&  .� \�E+   a��6   P'  � �   ��-  �-  Q'  � ^�E+  _� �   P'  \� �!   ��-  �-  Q'  � `'  �   W�-  S'  M� \E+   a�6   P+  ��     �.  -.  Q-+  � \.E+  a;�6   I   ;.  P.  Jh  �'  F:� $P.   	�#  P-.  w� @:   �p.  �.  Q;.  � QD.  �]]]r\z�6   Iq   �.  �.  Jh  M&  F:� -�.   	�#  P�.  �� �   ��.  �.  Q�.  � Q�.  �\�U.   I   �.  /  Jh  s&  F:� 2/   	�#  P�.  �� �   �4/  N/  Q�.  � Q/  �\�U.   I�   \/  q/  Jh  �&  F:� 7q/   	�#  PN/  �� �   ��/  �/  Q\/  � Qe/  �\�U.   I�   �/  �/  Jh  �&  F:� <�/   	�#  P�/  f� �   ��/  0  Q�/  � Q�/  �\�U.   I�   0  +0  Jh  @+  F:� A+0   	�#  P0  ��  :   �K0  o0  Q0  � Q0  �]]2\:�6   I   }0  �0  Jh  �&  F:� J�0   	�#  Po0  /� @   ��0  �0  Q}0  � Q�0  �\R00   I�   �0  �0  Jh  '  F:� O�0   	�#  P�0  �� `   �1  )1  Q�0  � Q�0  �\r00   I~   71  L1  Jh  1'  F:� TL1   	�#  P)1  f� �   �l1  �1  Q71  � Q@1  �\�00   bU  =�1   	;   b�   >�1  bB  ?�1  b�  E�1   	F   bB   F�1  bC  G�1  be  H�1  b8  I�1  b�  J�1  b

  X2   	Q   b�  Y2  b�
  Z2  c�   `12  	\   b�  fB2   	g   b�  gB2  b�  hB2  b�  nk2   	r   b�	  ok2  b�  pk2  bH  v�2   	}   b`  w�2  bw  x�2  b   y�2  b~  �2   	�   b   ��2  b�  ��2  b  ��2  b�   ��2  b�  ��2  b�	  ��2  b�  �"3   	�   b  �"3  b  �"3  b�  �"3  b�  �W3   	�   b�  �W3  b�  �W3  b�  �W3  bm  ��3   	�   b	  ��3  b2	  ��3  b�  ��3  b9  ��3  b[  ��3   	�   bJ  ��3  b�  ��3  b7  ��3  b�  �4   	�   bI	  �4  b$	  �4  b�   �+4   	�   bN  �+4  bp  �H4   	�   b�  �H4  b:  �H4  b�  �H4  bd   �H4  b�  ɉ4   	�   b  ʉ4  b�  ˉ4  b�	  Ѳ4   	�   b�  Ҳ4  b  ��4   	�   b�  ��4  b�  ��4  b�  ��4  b+  �5   	!  b�  �5  b�   �5  b  �-5   	!  b�
  �-5  b�  �-5  b  �V5   	!  b   �V5  bF  �V5  b�  �5   	"!  b�  �5  b�  �5  bD  O�5   	<!  b�  P�5  b1  Q�5  b�  W�5   	G!  b^  X�5  b�  3�5   	R!  b�  4�5  b�   86   	]!  b�  96  bl	  =(6  	h!  bN  >(6  b^  ?(6  bL  @(6  ba  D]6  	s!  bB  E]6  b�	  F]6  b  G]6  b  H]6  by  I]6  b�   �6   	~!  b�  !�6  �  �1  �6  :!   d>  Y  :!    6E   V9 �� �� �V  �I     4� std ) �)  v�/  w�/  {�/  �0  �40  �I0  �^0  ��0  ��0  ��0  ��0  �1  �;1  �[1  �|1  ��1  ��1  ��1  ��1  ��1  R2  U%2  [:2  \T2  b�2  cf4  eq4  f�4  g�4  h�4  i�4  j�4  k�4  l5  m65  qP5  ru5  t�5  u�5  v�5  x�5  y6  |6  ~'6  �96  �N6  �h6  �z6  ��6  ��6  ��6  ��6  5�6  68  768  @O8  %  0�=  �  �b  �3.  Fe  ��-  �3  �=  �  m8  s8   	�  
eq �<-  y8    s8  s8   
lt ��1  y8  :  s8  s8   ��  eF  �-  ^  �8  �8  �   �K  �9  �  x  �8   �(  
!  �8  �  �8  �  s8   1  �A  �8  �  �8  �8  �   �5  �'  �8  �  �8  �8  �   �3  �A  �8    �8  �  �   +  :  �  "  �8   	�  �C   �P  �  A  s8   �B  $6  y8  `  �8  �8   eof (�:  �  ?  ,N0  �  �8    _� ��-  �?  ��-  K  	\  �)   �e  	_�  �4  	c�8  �J  	d�8  ��  	q�  �  �8   ��  	s�    �8  �8   W  	y  �8  �-    	�  �J  
p�  �B  
k  �   %  
N/   �B  
Z  �8  N/  �8    �e  
y�  [V  
�  	k  �G  
!.   <  
x�  �4  
{�  �J  
|�  �J  
a+  `S  
��-  ~J  
��  �J  
��  �%  
�  �K  
�k   I  
�k  :!  
��8   %H  
��  �   �3  2�  �G  7/0  t3  B�8  �'  
��O  �8  V  
��N  y8  t  z  9   3  
�o+  y8  �  �  9   �P  
��O  �  �  �8   �M  
��P  �  �  �8   �,  
�-  �  �  �8  k   �+  
��R  N/  �    �8   3  
�   N/    +  �8  �8  �8   �/  !�B  �8  O  k  k  �8   �O  
�|6  b  m  �8  �8   (  ��6  �  �  �8  �8   �   
�-  N/  �  �  �8    �1  o�*  N/  �  �8  �8  k    �A  
$n%  N/  �  �  �8   �A  
(�I  N/      �8  N/   "A  
,�%  �8  (  .  �8   �1  
2E)  �  F  L  �8   �/  
6;&  �  d  j  �8   �>  
:�>  ~  �  �8   S  
A:2  k  �  �  �8  k  )0   �#  
K�(  �  �  �8  k  k  )0   9  
S>$  k  �  �  �8  k  k   -U  
[�7  y8       �8  )0   !�5  
d�-  @  N/  )0  k   !	1  
m�P  `  N/  )0  k   !�3  
v\-  �  N/  k  3.   !nU  
��-  �  N/  �  �   !nU  
�nG  �  N/  �  �   !nU  
��   �  N/  N/  N/   !nU  
�IP   	  N/  )0  )0   �J  
�rR  �-  	  k  k   �=  ��H  3	  H	  �8  k  k  k   V  �)  \	  b	  �8   "�'  
�D*  �8  #�0  
��	  �	  �8   $�0  ��	  �	  �8  �8   �0  ��	  �	  �8  �8   �0  ��	  �	  �8  �8  k  k   �0  ��	  
  �8  �8  k  k  �8   �0  �
  3
  �8  )0  k  �8   �0  �C
  S
  �8  )0  �8   �0  �c
  x
  �8  k  3.  �8   #�0  
"�
  �
  �8  �-   %�  
*,Q  �8  �
  �
  �8  �8   %�  
2�G  �8  �
  �
  �8  )0   %�  
=�%  �8  �
     �8  3.   %S� 
f�&  �      �8   %S� 
q�>  �  8  >  �8   &end 
y<  �  W  ]  �8   &end 
�6;  �  v  |  �8   %I 
��$  �  �  �  �8   %I 
��7  �  �  �  �8   %��  
�lC  �  �  �  �8   %��  
�CM  �  �  �  �8   %r 
��R  k      �8   %�K  
�r5  k  0  6  �8   %�3  
�j=  k  O  U  �8   '�� �  j  z  �8  k  3.   '�� 
��F  �  �  �8  k   %I  
v  k  �  �  �8   '�E  �|U  �  �  �8  k   '�1  
-�  �  �  �8   %�� 
5�?  y8      �8   %�:  
D�6  �  ,  7  �8  k   %�:  
UW  �  P  [  �8  k   &at 
k
/  �  s  ~  �8  k   &at 
��7  �  �  �  �8  k   %�F  
��/  �8  �  �  �8  �8   %�F  
�k:  �8  �  �  �8  )0   %�F  
��H  �8      �8  3.   %@  DA:  �8  &  1  �8  �8   %@  U�1  �8  J  _  �8  �8  k  k   %@  )�D  �8  x  �  �8  )0  k   %@  
��*  �8  �  �  �8  )0   %@  �6  �8  �  �  �8  k  3.   '�G  
-aN  �  �  �8  3.   (�3  �b*  �8      �8  �8   %�3  
^ 2  �8  1  F  �8  �8  k  k   %�3  �=  �8  _  o  �8  )0  k   %�3  
z�T  �8  �  �  �8  )0   %�3  
� @  �8  �  �  �8  k  3.   '� 
��E  �  �  �8  �  k  3.   %� 
�\+  �8  �    �8  k  �8   %� 
�u>  �8  (  B  �8  k  �8  k  k   %� g|=  �8  [  p  �8  k  )0  k   %� 
"�@  �8  �  �  �8  k  )0   %� 
9k<  �8  �  �  �8  k  k  3.   %� 
K�'  �  �  �  �8  �  3.   %bL  
d�R  �8  	    �8  k  k   %bL  
t�2  �  2  =  �8  �   %bL  �L&  �  V  f  �8  �  �   %�%  
�9F  �8    �  �8  k  k  �8   %�%  
�|<  �8  �  �  �8  k  k  �8  k  k   %�%  ��T  �8  �  �  �8  k  k  )0  k   %�%  
��A  �8    -  �8  k  k  )0   %�%  
b>  �8  F  `  �8  k  k  k  3.   %�%  
3%  �8  y  �  �8  �  �  �8   %�%  
'V7  �8  �  �  �8  �  �  )0  k   %�%  
<�+  �8  �  �  �8  �  �  )0   %�%  
Q'S  �8    "  �8  �  �  k  3.   %�%  
vj.  �8  ;  U  �8  �  �  N/  N/   %�%  
��9  �8  n  �  �8  �  �  )0  )0   %�%  
�C  �8  �  �  �8  �  �  �  �   %�%  
�>/  �8  �  �  �8  �  �  �  �   �?  ��&  �8       �8  k  k  k  3.   �1  �O  �8  8  R  �8  k  k  )0  k   ,)  
�z-  N/  v  k  3.  �8   )+E  �3J  N/  �  k  3.  �8   %�5  ��)  k  �  �  �8  N/  k  k   'n	 @D  �  �  �8  �8   %W�  
�6  )0       �8   %�A  
%�A  )0    %  �8   %��  
,Z5  �  >  D  �8   %�(  �;  k  ]  r  �8  )0  k  k   %�(  
I�%  k  �  �  �8  �8  k   %�(  
X�5  k  �  �  �8  )0  k   %�(  �^   k  �  �  �8  3.  k   %�(  
v�S  k      �8  �8  k   %�(  	K  k  /  D  �8  )0  k  k   %�(  
�o?  k  ]  m  �8  )0  k   %�(  J5  k  �  �  �8  3.  k   %NW  
��Q  k  �  �  �8  �8  k   %NW  /�I  k  �  �  �8  )0  k  k   %NW  
��,  k      �8  )0  k   %NW  
��;  k  /  ?  �8  3.  k   %�S  
��I  k  X  h  �8  �8  k   %�S  >T?  k  �  �  �8  )0  k  k   %�S  
05  k  �  �  �8  )0  k   %�S  
$S:  k  �  �  �8  3.  k   %�>  
2hL  k      �8  �8  k   %�>  SUB  k  *  ?  �8  )0  k  k   %�>  
Q�2  k  X  h  �8  )0  k   %�>  _�K  k  �  �  �8  3.  k   %�4  
qT  k  �  �  �8  �8  k   %�4  j�K  k  �  �  �8  )0  k  k   %�4  
��5  k      �8  )0  k   %�4  N.  k  *  :  �8  3.  k   %U+  
�)  "  S  c  �8  k  k   %��  
�!1  �-  |  �  �8  �8   %��  ��T  �-  �  �  �8  k  k  �8   %��  ��O  �-  �  �  �8  k  k  �8  k  k   %��  �;.  �-      �8  )0   %��  ��B  �-  *  ?  �8  k  k  )0   %��  ��,  �-  X  r  �8  k  k  )0  k   	  *!T  3.  +�E  �  +�F  �   ,�&  ,�7  	"  �o  >�   �| C�-  -Q  b�   	�  -�F c�  -�R  d�  -3  e�  -�  f�  -�K  g�  -�@  h�   .all i�  ?/�� �}  :!  ��8   NF  �F9  �E  ��  p0  �F9  �%  ��1  0S  �R9  0�R  �R9  03  �R9  0�$  �R9  0�K  �R9  0�@  �R9  0�@  �]9  �4  �Z  �  �  9   �=  y)  �  �  9   1��     9  s9  �   1�� .  >  9  )0  �   1�� N  Y  9  �   1N  i  t  9  �-   1�� �  �  9  s9   �  �U  �  �  9  s9   �&  �.  y8  �  �  9   �F  &�;  �  �  9  y9  �   �9  )�Q      9  y9  h9   WR  ,`2  (  8  9  y9  @9   �S  /=  L  \  9  @9  L9   2e  7,  l  9  L9  �    �$  9   0OD  9  0gP  9  0�F  $9  3< #  4��  ґr  �  e>  )0  A)   4�h  �ܧ  �  e>   5��  ��  A)    e>   6�< �; A)  A)  )0    7id ��  �U  ��   0�I  ��8  �  �<?  ]  h  49  :9   8id �w  �  49  :9   9id ��  �  49   :4H  ��(  �  �  @9    �o  u�  �  "9   �o  ~�  �  "9  (9   $�o  ��     "9  )0   �o  �  %  "9  (9  )0  �   �o  �5  J  "9  (9  (9  �   5  �Z  e  "9  �-   (�  ��*  (9  }  �  "9  (9   (H�  ��N  �   �  �  .9   (U  �9  y8  �  �  .9  (9   (2  �t*  y8  �  �  .9  (9   ;jP  �D  �     (9   <RD  �Q  (9  =�o  7(   3   "9  9   >�K  :�N  >�A  =�5  �K  @I  �  e   �   �,  CH<  y   �   "9  (9  (9  �   	#  	�  	'   	�  � >"  ?W  3=!  @�4  @�$  @q-  @c=  @o'  @�5   @�%  � @�8  �@X)  �@�%  �@�  �@aO  �@Y=  � @P  �� @�C  ��@wS  �@�O  � @�?  �@�5  �� ?
$ gv!  @)W  @�   @�U  @�A  @�8  @�P   @EH  �� ?�4  ��!  @O   @�7  @(  @�Q  @G  �� 3b4 +#  A�  Jv!  �P  ��   B�4  �!  	�!  Cdec �!  Bt-  �!  Chex �!  Br'  �!  B< �!   Coct �!  @B� �!  �D[)  �!   D�%  "�!   D�  &�!   DdO  )�!   D\=  ,�!   D�P  /�!    D�C  3�!   @BzS  6�!  �B�O  9�!  JD�?  <�!  B(  Q�"  	�!  B�Q  V�"  BO  Y�"   A�9  i=!  Cin w#  	�"  Cout z#   <�9  =9  >�9  @%:  A0:  BJ:  Ce:  D�:  E�:  F�:  G�:  H�:  ד  ��#  ��  ��  � �N/  �4  ��8  *{�  N/   ?�0 ��#  @R1 @�1  @�1 @�2 @�3  ?F2 � $  @/ @v/  @�4  	�#  	�#  |� �%  E�+ �8  E}�   �8  E�. !�8  E�3 &�8  E�. '�8   EJ- (�8   E_5 )�8  F�4 1�8  �Fr6 2�8  [Ef1 3�8  �E0 4�8  &E/, 6�8  E�1 7�8  EY2 8�8  EV, 9 $  E5 ;�8   Ex, J�8  E�+ L�8  E�2 M�8   E�4 O�8   E�3 P�8   E�0 R$  min �� �-  max �� �-  "T4 ,Y� �-  "/5 / � �-  "�2 ?0� �-  "�1 B�� �-  "]2 E�� �-  "�4 H^� �-   �� \g'  E�+ ^�8  E}�  k�8  5E�. l�8  E�3 q�8  E�. r�8   EJ- s�8   E_5 t�8  F�4 |�8  �xFr6 }�8  �}Gf1 ~�8   G0 �8  4E/, ��8  E�1 ��8  EY2 ��8  EV, � $  E5 ��8   Ex, ��8  E�+ ��8  E�2 ��8   E�4 ��8   E�3 ��8   E�0 �$  min ap� �-  max d� �-  "T4 w�� �-  "/5 z�� �-  "�2 �� �-  "�1 �9� �-  "]2 �T� �-  "�4 ��� �-   �� �)  E�+ ��8  E}�  ��8  @E�. ��8  E�3 ��8  E�. ��8   EJ- ��8   E_5 ��8  F�4 ��8  ��Fr6 ��8  �YGf1 ��8   @G0 ��8  DE/, ��8  E�1 ��8  EY2 ��8  EV, � $  E5 ��8   Ex, ��8  E�+ ��8  E�2 ��8   E�4 ��8   E�3 ��8   E�0 �$  min ��� �-  max �/� �-  "T4 ��� �-  "/5 �H� �-  "�2 �� �-  "�1 ��� �-  "]2 �~� �-  "�4 ��� �-   h�  1!o  <)  )0  U;  [;  a;   	A)  W�  1g;  	�  <�  r��  u)  )0  p<  [;  a;   �  ��l  �)  )0  j=  [;  a;   H�8 R#< )0    I$   %E�-  �  $,�  -�  K  :\+  �e  =�  � ?N/  "  @)0  �4  A�8  �J  B�8  �A  O#*  )*  �8   �A  Q9*  D*  �8  �8   �A  VT*  _*  �8  �-   (�
 Y51  �)  w*  �*  �8  �)   (�
 ]�R  �)  �*  �*  �8  *   (� c?  �)  �*  �*  �8  �)  �0   J_ m.   �*  �*  �8  �)  �)   (�3  q89  �)  	+  +  �8   J.E  ��3  #+  3+  �8  �)  �8   J�(  ��(  G+  R+  �8  �)   K_Tp 3.   	�)  LZD  ��-  MF�  �N/   A��  ��#  A�4  ��#  A� ��#  #��  ��+  �+  ;   N��  ��+  �+  ;  ;   %*  ��}  �+  �+  �+  ;   %Ư  �?s  �+  ,  ,  ;   %�F  �Ϭ  %;  -,  3,  ;   %�F  ��  a+  L,  W,  ;  �-   %a�  �
�  %;  p,  v,  ;   %a�   ��  a+  �,  �,  ;  �-   %�:  ,�  �+  �,  �,  ;  |+   %�F  		n  %;  �,  �,  ;  |+   %(*  ��  a+  �,  -  ;  |+   % I  h�  %;  -  *-  ;  |+   %�O  7k  a+  C-  N-  ;  |+   %WC  ]�  ;  g-  m-  ;   *{�  N/  *�  "   ,8E  	a+  O�� �cD   P�  Po  P�  P�  P�  P�  P�	  Qint P(  P#  P�� P�� P�� _� ԫ-  �  �-  pW   �-  qW  !�-    "�-    #�-  P�  Rs  N�-  �  V�-  SFd .  .  <.  `  D�-  �  W.  �  _.  �  e�-  t   m�-  a  u�-    ~�-  �  ��-  3  ��-  �  ��-  H  ��-  y  ��-    ��-  s  ��-  T   ��-  �  ��-  F  ��-  �  ��-  �  ��-    ��-  V  ��-  T3.  P�  \	  2�-  o  7�-  �  <�-  �  C�-  �  �-  T�-  U*  �/  �  �-   Vrem �-   +   �/  U#@  �/  �  $�-   Vrem %�-   A  &�/  W� ��-  0  0   T0  XW�  >�-  )0  )0   T/0  	3.  W�  H�-  I0  )0   W�  I�-  ^0  )0   W�  �:.  �0  �0  �0  �-  �-  �0   T�0  YT�0  Z�-  �0  �0  �0   [div �/  �0  �-  �-   W    �N/  �0  )0   \�   �/  �0  �-  �-   \�  .�-  1  )0  �-   \�  \�-  .1  .1  )0  �-   T41  P  \3  >�-  [1  .1  )0  �-   ]�  |1  :.  �-  �-  �0   ^k� q�-  _�  |�1  �-   W  W�-  �1  )0  �1   TN/  W  f�-  �1  )0  �1  �-   W�  g�-  �1  )0  �1  �-   W?  ��-  2  )0   W��  E�-  %2  )0  )0   W��  UN/  :2  �-   W��  ON/  T2  N/  )0   W��  F�-  s2  N/  )0  �-   	\   (.  gX   (.  X\  !&�2  X\  X!,�3  $Z  !.R.   \ !/�-  � !1�/  Z  !2�-  K]  !3�-  �_  !4�-  \W  !5�-  �Z  !6�-  -_  !8�3   VY  !9�3  $`  !:4  (�Y  !;4  ,7_  !<04  0BY  !=O4  4b\  !>04  8\  !?04  <7Y  !@04  @ Z  !A`4  DSX  !B`4  Hn4 !D.  L`  !F�3  P*5 !G�3  T Z~2  �3  :.  �-  �3   T�2  T�3  Z~2  �3  �0  �-  �3   T�3  Z�-  4  �3  s2  �-   T�3  Zs2  4  �3   T4  Z�-  04  �3   T!4  Z�3  O4  )0  )0  �3   T64  ``4  �3   TU4  �^  "!s2  ]Z  "1�4  �4   T�2  WaY  "��-  �4  �4   \\  "C�-  �4  �4   \xZ  "M�-  �4  �4   W`  "��-  �4  �4   \�^  "r�-  �4  �4   \_X  "��-  5  �4  5   Tf4  \�_  "�N/  65  N/  �-  �4   W�\  "��4  P5  )0  )0   \4Z  "��-  u5  �0  �-  �-  �4   W7`  "��4  �5  )0  )0  �4   \>]  "	�-  �5  �4  �-  �-   \�Z  "�-  �5  �4  �5   T�5  	f4  \�Y  " �-  �5  �4   \�Y  "��-  6  �4   a\  "��-  W�_  0N/  '6  N/   ]�]  "W96  )0   WD[  "T�-  N6  )0   W�[  "a�-  h6  )0  )0   ]�\  ")z6  �4   _Y@ "��6  �4  N/   W�[  "��-  �6  �4  N/  �-  �-   ^�]  "i�4  WD]  "wN/  �6  N/   \}W  "��-  �6  �-  �4   �  8#8  �{  #N/   ]�  #N/  \�  # N/  �D  #!N/  �3  #"N/  U>  ##N/  &�  #$N/  �  #%N/  �*  #&N/   ڡ  #'3.  $�U  #(3.  %TL  #)3.  &�I  #*3.  'Q  #+3.  (�C  #,3.  )�J  #-3.  *1  #.N/  ,o(  #/3.  0�U  #03.  1PL  #13.  2�I  #23.  3Q  #33.  4�C  #43.  5�J  #53.  6 W)%  #KN/  68  �-  )0   ^GT  #PA8  T�6  b$pO qO $!G8  I2*  7m8  c8�   d�  d�  P�  T�  T�  d"  d3.  d/0  T�)  d\+  T\+  T�  d  �  & �-  	�-  	y8  T.  T�  T"  T  d  d�  d"  e�-  9  f Tr  T'  	9  T9  	)0  T�  d�   T�   T#  d�   T�   TL9  T�   e@9  ]9  f eh9  h9  f Tn9  	@9  d�   T�   �l  '�-  j�  '#�-  gtm ,',%:  ,g  '.�-   �  '/�-  �  '0�-  ��  '1�-  ��  '2�-  ��  '3�-  ��  '4�-  �  '5�-  d�  '6�-   ��  '7�-  $~�  '8)0  ( ^\�  '>�9  Wѯ  'H�-  J:  9  9   W��  'M9  _:  _:   T�9  W�  'C9  z:  z:   T9  W#�  'aN/  �:  �:   T�:  	�9  W�� 'fN/  �:  �:   T�:  	9  W��  'W_:  �:  �:   W[v  '\_:  �:  �:   W��  'R�-  ;  N/  �-  )0  �:   Ta+  d;  	N/  T�-  da+  hv%  hF%  h&'  h�&  h`  h�(  h�(  d�-  d�!  d<)  T�-  i)  �  �a<  j__s 1)0  � j__v 1a<  �k�*  1f<  �lk<  �m8I N<  n'U  5N/  l� nR'  6L)  �� ngw  7N/  �� o�� :N/  �\nN� ;y8  �� p�8  p��D  p��D  p��D  p�8  p��D  pK8  pS�D   p��D  p�E   	U;  	[;  	a;  d�-  iQ)  �$  �[=  j__s r)0  � j__v r[=  �k�*  r`=  �le=  �mPI H=  n'U  vN/  �� nR'  wL)  � ngw  xN/  ,� o�� {N/  �\p�8  p��D  p��D  p��D  p8  p�1  pk8  ps�D   p��D  p�E   	p<  	[;  	a;  d�-  iu)  �  �V>  j__s �)0  � j__v �V>  �k�*  �[>  �l`>  �mhI C>  n'U  �N/  U� nR'  �L)  ~� ngw  �N/  �� q__p ��-  �� p8  p�D  p&�D  p4�D  pB8  pS!E  p�8  r��D   p��D  pE   	j=  	[;  	a;  dA)  i�  4   ��>  k(�  ҭ>  � s__s �)0  � lA)  �pD�)   	e>  i�  P   ��>  k(�  ��>  �  	e>  i�  `   ��>  l�>  �  	e>  i  p   �?  lA)  � l)0  � tD  O*?   	<.  t�  P*?  t1  Q*?  t�  WS?   	G.  t^  XS?  tU  =p?   	\.  t�   >p?  tB  ?p?  t�  E�?   	g.  tB   F�?  tC  G�?  te  H�?  t8  I�?  t�  J�?  t

  X�?   	r.  t�  Y�?  t�
  Z�?  u�   `@  	}.  t�  f @   	�.  t�  g @  t�  h @  t�  nI@   	�.  t�	  oI@  t�  pI@  tH  vr@   	�.  t`  wr@  tw  xr@  t   yr@  t~  �@   	�.  t   ��@  t�  ��@  t  ��@  t�   ��@  t�  ��@  t�	  ��@  t�  � A   	�.  t  � A  t  � A  t�  � A  t�  �5A   	�.  t�  �5A  t�  �5A  t�  �5A  tm  �jA   	�.  t	  �jA  t2	  �jA  t�  �jA  t9  �jA  t[  ��A   	�.  tJ  ��A  t�  ��A  t7  ��A  t�  ��A   	�.  tI	  ��A  t$	  ��A  t�   �	B   	�.  tN  �	B  tp  �&B   	�.  t�  �&B  t:  �&B  t�  �&B  td   �&B  t�  �gB   	/  t  �gB  t�  �gB  t�	  ѐB   	/  t�  ҐB  t  حB   	/  t�  ٭B  t�  ڭB  t�  ۭB  t+  ��B   	"/  t�  ��B  t�   ��B  t  �C   	-/  t�
  �C  t�  �C  t  �4C   	8/  t   �4C  tF  �4C  t�  �]C   	C/  t�  �]C  t�  �]C  t�  3�C   	[/  t�  4�C  t�   8�C   	f/  t�  9�C  tl	  =�C  	q/  tN  >�C  t^  ?�C  tL  @�C  ta  D�C  	|/  tB  E�C  t�	  F�C  t  G�C  t  H�C  ty  I�C  t�   BD   	�/  t�  !BD  e)0  cD  vT/   	SD  w�-  �	x�  �� �	WY2  Q�-  �D  )0   )�  (��  :.  �D  �   y�d  :.  �D  :.  �0  T/   W�� V�-  �D  )0  �1   �e  (�Ӫ  �D  :.   z>  Y  E  :.   {  !E  :.   |� "D�-  )0  )0  }  C5   A ^� �� �V  �I     �� (  _� �7   �  �  8k  �{  k   ]�  k  \�   k  �D  !k  �3  "k  U>  #k  &�  $k  �  %k  �*  &k   ڡ  'q  $�U  (q  %TL  )q  &�I  *q  'Q  +q  (�C  ,q  )�J  -q  *1  .k  ,o(  /q  0�U  0q  1PL  1q  2�I  2q  3Q  3q  4�C  4q  5�J  5q  6 q  �  std # "  5>   6"  7D"  @�#  	%  0�=  �n  �b  �q  Fe  �2"  
�3  �=  �  (  (   �  eq �<-  (    (  (   lt ��1  (  !  (  (   ��  eF  2"  E  $(  $(  n   �K  �9  n  _  $(   �(  
!  $(  �  $(  n  (   1  �A  *(  �  *(  $(  n   �5  �'  *(  �  *(  $(  n   �3  �A  *(  �  *(  n  �   +  :  �  	  0(   �  �C   �P  �  (  (   �B  $6  (  G  0(  0(   eof (�:  �  ?  ,N0  �  0(    _� 	�7   �?  	�%   K  
\  )$   �e  
_n  �4  
c6(  �J  
d<(  ��  
q�  �  T(   ��  
s�  �  T(  Z(   W  
y�  T(  2"    �  �J  pz  �B  R  �   %  k   �B  A  x(  k  Z(    �e  y�  [V  k  R  �G  !   <  x�  �4  {�  �J  |�  �J  �%  `S  ��'  ~J  �z  �J  �  �%  �  �K  �R   I  �R  :!  �m(   %H  ��  �   �3  2k  �G  7?"  t3  B�(  �'  ��O  �(  V  ��N  (  [  a  �(   3  �o+  (  x  ~  �(   �P  ��O  �  �  �(   �M  ��P  �  �  �(   �,  �-  �  �  �(  R   �+  ��R  k  �  �  �(   3  �   k      �(  Z(  Z(   �/  !�B  �(  6  R  R  Z(   �O  �|6  I  T  �(  Z(    (  ��6  h  s  �(  Z(   !�   �-  k  �  �  �(   "�1  o�*  k  �  �(  Z(  R    !�A  $n%  k  �  �  ~(   !�A  (�I  k  �  �  �(  k   !"A  ,�%  �(      ~(   !�1  2E)  �  -  3  ~(   !�/  6;&  �  K  Q  ~(    �>  :�>  e  k  �(   !S  A:2  R  �  �  ~(  R  9"    �#  K�(  �  �  ~(  R  R  9"   !9  S>$  R  �  �  ~(  R  R   !-U  [�7  (  �    ~(  9"   #�5  d�-  '  k  9"  R   #	1  m�P  G  k  9"  R   #�3  v\-  g  k  R  q   #nU  ��-  �  k  �  �   #nU  �nG  �  k  �  �   #nU  ��   �  k  k  k   #nU  �IP  �  k  9"  9"   �J  �rR  2"  	  R  R    �=  ��H  	  /	  �(  R  R  R    V  �)  C	  I	  �(   $�'  �D*  �(  %�0  �j	  p	  �(   &�0  ��	  �	  �(  Z(   �0  ��	  �	  �(  �(   �0  ��	  �	  �(  �(  R  R   �0  ��	  �	  �(  �(  R  R  Z(   �0  �
  
  �(  9"  R  Z(   �0  �*
  :
  �(  9"  Z(   �0  �J
  _
  �(  R  q  Z(   %�0  "p
  {
  �(  2"   '�  *,Q  �(  �
  �
  �(  �(   '�  2�G  �(  �
  �
  �(  9"   '�  =�%  �(  �
  �
  �(  q   'S� f�&  �       �(   'S� q�>  �    %  ~(   (end y<  �  >  D  �(   (end �6;  �  ]  c  ~(   'I ��$  �  |  �  �(   'I ��7  �  �  �  ~(   '��  �lC  �  �  �  �(   '��  �CM  �  �  �  ~(   'r ��R  R  �  �  ~(   '�K  �r5  R      ~(   '�3  �j=  R  6  <  ~(   )�� �  Q  a  �(  R  q   )�� ��F  v  �  �(  R   'I  v  R  �  �  ~(   )�E  �|U  �  �  �(  R   )�1  -�  �  �  �(   '�� 5�?  (  �  �  ~(   '�:  D�6  �      ~(  R   '�:  UW  �  7  B  �(  R   (at k
/  �  Z  e  ~(  R   (at ��7  �  }  �  �(  R   '�F  ��/  �(  �  �  �(  �(   '�F  �k:  �(  �  �  �(  9"   '�F  ��H  �(  �  �  �(  q   '@  DA:  �(      �(  �(   '@  U�1  �(  1  F  �(  �(  R  R   '@  )�D  �(  _  o  �(  9"  R   '@  ��*  �(  �  �  �(  9"   '@  �6  �(  �  �  �(  R  q   )�G  -aN  �  �  �(  q   *�3  �b*  �(  �  �  �(  �(   '�3  ^ 2  �(    -  �(  �(  R  R   '�3  �=  �(  F  V  �(  9"  R   '�3  z�T  �(  o  z  �(  9"   '�3  � @  �(  �  �  �(  R  q   )� ��E  �  �  �(  �  R  q   '� �\+  �(  �  �  �(  R  �(   '� �u>  �(    )  �(  R  �(  R  R   '� g|=  �(  B  W  �(  R  9"  R   '� "�@  �(  p  �  �(  R  9"   '� 9k<  �(  �  �  �(  R  R  q   '� K�'  �  �  �  �(  �  q   'bL  d�R  �(  �     �(  R  R   'bL  t�2  �    $  �(  �   'bL  �L&  �  =  M  �(  �  �   '�%  �9F  �(  f  {  �(  R  R  �(   '�%  �|<  �(  �  �  �(  R  R  �(  R  R   '�%  ��T  �(  �  �  �(  R  R  9"  R   '�%  ��A  �(  �    �(  R  R  9"   '�%  b>  �(  -  G  �(  R  R  R  q   '�%  3%  �(  `  u  �(  �  �  �(   '�%  'V7  �(  �  �  �(  �  �  9"  R   '�%  <�+  �(  �  �  �(  �  �  9"   '�%  Q'S  �(  �  	  �(  �  �  R  q   '�%  vj.  �(  "  <  �(  �  �  k  k   '�%  ��9  �(  U  o  �(  �  �  9"  9"   '�%  �C  �(  �  �  �(  �  �  �  �   '�%  �>/  �(  �  �  �(  �  �  �  �   !�?  ��&  �(  �    �(  R  R  R  q   !�1  �O  �(    9  �(  R  R  9"  R   ,)  �z-  k  ]  R  q  Z(   ++E  �3J  k  �  R  q  Z(   '�5  ��)  R  �  �  ~(  k  R  R   )n	 @D  �  �  �(  �(   'W�  �6  9"  �  �  ~(   '�A  %�A  9"      ~(   '��  ,Z5  }  %  +  ~(   '�(  �;  R  D  Y  ~(  9"  R  R   '�(  I�%  R  r  �  ~(  �(  R   '�(  X�5  R  �  �  ~(  9"  R   '�(  �^   R  �  �  ~(  q  R   '�(  v�S  R  �  �  ~(  �(  R   '�(  	K  R    +  ~(  9"  R  R   '�(  �o?  R  D  T  ~(  9"  R   '�(  J5  R  m  }  ~(  q  R   'NW  ��Q  R  �  �  ~(  �(  R   'NW  /�I  R  �  �  ~(  9"  R  R   'NW  ��,  R  �  �  ~(  9"  R   'NW  ��;  R    &  ~(  q  R   '�S  ��I  R  ?  O  ~(  �(  R   '�S  >T?  R  h  }  ~(  9"  R  R   '�S  05  R  �  �  ~(  9"  R   '�S  $S:  R  �  �  ~(  q  R   '�>  2hL  R  �  �  ~(  �(  R   '�>  SUB  R    &  ~(  9"  R  R   '�>  Q�2  R  ?  O  ~(  9"  R   '�>  _�K  R  h  x  ~(  q  R   '�4  qT  R  �  �  ~(  �(  R   '�4  j�K  R  �  �  ~(  9"  R  R   '�4  ��5  R  �  �  ~(  9"  R   '�4  N.  R    !  ~(  q  R   'U+  �)  	  :  J  ~(  R  R   '��  �!1  2"  c  n  ~(  �(   '��  ��T  2"  �  �  ~(  R  R  �(   '��  ��O  2"  �  �  ~(  R  R  �(  R  R   '��  �;.  2"  �  �  ~(  9"   '��  ��B  2"    &  ~(  R  R  9"   '��  ��,  2"  ?  Y  ~(  R  R  9"  R     ,!T  q  -�E  �  -�F  �   .�&  .�7  	  �o  >2   �| C2"  /Q  b�   �  /�F c�  /�R  d�  /3  e�  /�  f�  /�K  g�  /�@  h�   0all i�  ?1�� �d  :!  �m(   NF  ��(  �E  �n  p0  ��(  �%  ��(  2S  ��(  2�R  ��(  23  ��(  2�$  ��(  2�K  ��(  2�@  ��(  2�@  �
)   �4  �Z  �  �  �(    �=  y)  �  �  �(   3�� �    �(   )  n   3��   %  �(  9"  n   3�� 5  @  �(  n   3N  P  [  �(  2"   3�� k  v  �(   )    �  �U  �  �  �(   )   !�&  �.  (  �  �  �(    �F  &�;  �  �  �(  &)  �    �9  )�Q  �  �  �(  &)  )    WR  ,`2      �(  &)  �(    �S  /=  3  C  �(  �(  �(   4e  7,  S  �(  �(  n    �$  �(   2OD  �(  2gP  �(  2�F  $�(  5< �  6< r�  �-  n    7id �H  �U  �n   2�I  �m(   �  �<?  �  �  �(  �(   8id �    �(  �(   9id �&  ,  �(   :4H  ��(  n  A  �(    �o  uX  ^  �(   �o  ~n  y  �(  �(   &�o  ��  �  �(  9"   �o  ��  �  �(  �(  9"  �   �o  ��  �  �(  �(  �(  �   5  ��  �  �(  2"   *�  ��*  �(      �(  �(   *H�  ��N  7   4  :  �(   *U  �9  (  R  ]  �(  �(   *2  �t*  (  u  �  �(  �(   ;jP  �D  �  �  �(   <RD  �Q  �(  =�o  7�  �  �(  �(   >�K  :�N  >�A  =�5  �K  @I  �  �  �    �,  CH<     "   �(  �(  �(  �   �  �     �  � >	  <7)  =,)  >B)  @�)  A�)  B�)  C*  D-*  EM*  Fm*  G�*  H�*  ד  ��   ��  �y  � �k  �4  �6(  ,{�  k   v�*  w-+  {8+  �T+  �i+  �~+  ��+  ��+  ��+  �,  �!,  �<,  �\,  �|,  ��,  ��,  ��,  ��,  ��,  �-  R&-  U@-  [U-  \o-  5��  �!  ?�E  *e�  �!  �!  �-  k  n  9"  B*   ?ƙ  =��  �!  �!  �.  "   ,!T  q   u!  n  @�  "  A�  z�!  "  �.  n   ,!T  q   W�  1�.   B)%  Kk  2"  2"  9"   Cint ?"  q  DGT  PO"  >   �  `"  �  �  o  �	  �  qW  !2"    "�"  �  #  .  <�"  `  D2"  �  W�"  �  _�"  �  e2"  t   m2"  a  u2"    ~2"  �  �2"  3  �2"  �  �2"  H  �2"  y  �2"    �2"  s  �2"  T   �2"  �  �2"  F  �2"  �  �2"  �  �2"    �2"  V  �2"  �  Es  NU"  �  VU"  \	  22"  o  72"  �  <2"  �  C2"  �  2"  �#  FGpO qO !�#  H$   E�'  	�  $,n  -y  K  :�%  �e  =n  � ?k  "  @9"  �4  A6(  �J  B<(  �A  O�$  �$  B(   �A  Q�$  �$  B(  H(   �A  V�$  �$  B(  2"   *�
 Y51  A$  �$  �$  N(  Y$   *�
 ]�R  M$  �$  %  N(  e$   *� c?  A$  %  +%  B(  5$  �#   ?_ m.   ?%  O%  B(  A$  5$   *�3  q89  5$  g%  m%  N(   ?.E  ��3  �%  �%  B(  A$  <(   ?�(  ��(  �%  �%  B(  A$   I_Tp q   )$  JZD  ��'  KF�  �k   L��  ��   L�4  ��   L� ��   %��  �&  &  �*   M��  �)&  4&  �*  �*   '*  ��}  �%  M&  S&  �*   'Ư  �?s  �%  l&  r&  �*   '�F  �Ϭ  �*  �&  �&  �*   '�F  ��  �%  �&  �&  �*  2"   'a�  �
�  �*  �&  �&  �*   'a�   ��  �%  �&  �&  �*  2"   '�:  ,�  �%  '  '  �*  �%   '�F  		n  �*  5'  @'  �*  �%   '(*  ��  �%  Y'  d'  �*  �%   ' I  h�  �*  }'  �'  �*  �%   '�O  7k  �%  �'  �'  �*  �%   'WC  ]�  �*  �'  �'  �*   ,{�  k  ,�  	   .8E  �%   �� �� �� H2*  7(  N8�   O�  O�  �  �  �  O	  Oq  O?"  )$  O�%  �%  �  O  f(    �   2"    �  	    O  O�  O	  P7   �(  Q Y    �(  �(  9"  �  O2   2   �  O"   "   �(  '   k  P�(  
)  Q P)  )  Q )  �(  O,   ,   �l  %   j�  #%   Rtm ,,�)  ,g  .2"   �  /2"  �  02"  ��  12"  ��  22"  ��  32"  ��  42"  �  52"  d�  62"   ��  7%   $~�  89"  ( D\�  >7)  Bѯ  H�'  �)  ,)  ,)   B��  M,)  *  *   B)  B�  C,)  '*  '*   ,)  B#�  ak  B*  B*   H*  B)  B�� fk  b*  b*   h*  ,)  B��  W*  �*  b*   B[v  \*  �*  b*   B��  R,   �*  k  ,   9"  B*   �%  O�*  k  �'  O�%  S *  �*  �   2"   Trem  2"   +    �*  S #@  -+  �   $%    Trem  %%    A   &+  B�  �2"  M+  M+   S+  UB�   >�'  i+  9"   B�   H2"  ~+  9"   B�   I%   �+  9"   B�   �#  �+  �#  �#  ,   ,   �+   �+  V2"  �+  �#  �#   Wdiv  �*  �+  2"  2"   B     �k  ,  9"   X�    -+  !,  %   %    X�   .2"  <,  9"  ,    X�   \,   \,  `(  9"  ,    X3   >2"  |,  `(  9"  ,    Y�   �,  �#  ,   ,   �+   Dk�  q2"  Z�   |�,  |"   B   W�'  �,  9"  �(   B   f%   �,  9"  �(  2"   B�   g7   -  9"  �(  2"   B?   �2"  &-  9"   B��  !E2"  @-  9"  9"   B��  !Uk  U-  2"   B��  !Ok  o-  k  9"   B��  !F,   �-  k  9"  ,    �  [�  �-  �-  \h  �-  ]4&  rn   �-  �!  ^~!  ��   ��-  �.  _h  �.  � `__s +k  �aǆ  +n  �a�l  +9"  �ay  ,B*  �b�n   �.  c'U  .k  .� c�� /�!  L� cgw  0k  _� cR'  3�!  s� d�"  d��4  d��4  d��4  d�"  d��*  d�"  d��4   d5  d"5   �-  �!  [�!  �.  �.  \h  �.  e4&  zn   �.  u!  2"  ^�!   H  �/  u/  _h  u/  � f"  �g�.  ��  Ak/  h�.   i�.  Pj�-  �   �h�-   i�-  P  d�15   �.  kU  =�/   �"  k�   >�/  kB  ?�/  k�  E�/   �"  kB   F�/  kC  G�/  ke  H�/  k8  I�/  k�  J�/  k

  X�/   �"  k�  Y�/  k�
  Z�/  l�   `%0  �"  k�  f60   �"  k�  g60  k�  h60  k�  n_0   �"  k�	  o_0  k�  p_0  kH  v�0   �"  k`  w�0  kw  x�0  k   y�0  k~  �0   �"  k   ��0  k�  ��0  k  ��0  k�   ��0  k�  ��0  k�	  ��0  k�  �1   �"  k  �1  k  �1  k�  �1  k�  �K1   
#  k�  �K1  k�  �K1  k�  �K1  km  ��1   #  k	  ��1  k2	  ��1  k�  ��1  k9  ��1  k[  ��1    #  kJ  ��1  k�  ��1  k7  ��1  k�  ��1   +#  kI	  ��1  k$	  ��1  k�   �2   6#  kN  �2  kp  �<2   A#  k�  �<2  k:  �<2  k�  �<2  kd   �<2  k�  �}2   L#  k  �}2  k�  �}2  k�	  Ѧ2   W#  k�  Ҧ2  k  ��2   b#  k�  ��2  k�  ��2  k�  ��2  k+  ��2   m#  k�  ��2  k�   ��2  k  �!3   x#  k�
  �!3  k�  �!3  k  �J3   �#  k   �J3  kF  �J3  k�  �s3   �#  k�  �s3  k�  �s3  kD  O�3   �#  k�  P�3  k1  Q�3  k�  W�3   �#  k^  X�3  k�  3�3   �#  k�  4�3  k�   8�3   �#  k�  9�3  kl	  =4  �#  kN  >4  k^  ?4  kL  @4  ka  DQ4  �#  kB  EQ4  k�	  FQ4  k  GQ4  k  HQ4  ky  IQ4  k�   �4   �#  k�  !�4  BY2  !Q,   �4  9"   +�  "��  �#  �4  n   m�d  �#  �4  �#  �#  �#   
�e  "�Ӫ  5  �#   n>  Y  "5  �#   o  15  �#   p�  "��  �#  n    �   �G � �� �b �I     �� std  �  v  6�  x  K�  �  M�   x  Ob   m   �  �   	�  Qw  �   �   �   	�  R  �   �   �   
  T8  �  �   �   �   x  Z�   �   �   x  \�   �   �  �   x  _�     �  �   x  c  #  �  �   �  p�  �  ;  F  �  �   �  t�  �  ^  i  �  �   �  {y  �  �  �   n	 ~%  �  �  �  �   �  ��  �  �  �  �   �  �h  �  �  �    ;    :;   �  ��  � �  �S L%  0@!  _� ��  0�  1�  2�  3�  5>  6T  7j  8�  :�  ;�  <  =(  ?�  @�  B�  C�  D�  E�  GI  H_  Iu  J�  L�  M  N  O3  Q�  R�  �?  �0  5A  6n  7�  � 	'��  
)� ��  �  �   � :  @  �   �� �  V  a  �  �   (� "�     }  �    ��   	[ O�   �  6y 	)�     Ic  
1�      ;   �   �  !�  ";    ;   #int $�  �  $�  $�  $o  $�  $�  $�  $�	  $(  $#  $   �_  �  $,  -�   $�� $�� $�� 2*  7�  %8   $�  �    �  "  �O   �O )  pW     qW  !�    "    #7  ` &"  ` '  �^ ()  �^ )  �T *�  �T +  iY ,7  hY -  �e 0"  �e 1  [ 2�  [ 3  Q 4�  Q 5  �_ 67  �_ 7  �] :�  �] ;  �Q >7  �Q ?  .  <�  `  D�  �  W�  �  _�  �  e�  t   m�  a  u�    ~�  �  ��  3  ��  �  ��  H  ��  y  ��    ��  s  ��  T   ��  �  ��  F  ��  �  ��  �  ��    ��  V  ��  �  $�  s  N�  �  V�  \	  2�  o  7�  �  <�  �  C�  �  �    �  &pO qO !  $Ye $�[ $  '�  8n  �{  �   ]�  �  \�   �  �D  !�  �3  "�  U>  #�  &�  $�  �  %�  �*  &�   ڡ  '�  $�U  (�  %TL  )�  &�I  *�  'Q  +�  (�C  ,�  )�J  -�  *1  .�  ,o(  /�  0�U  0�  1PL  1�  2�I  2�  3Q  3�  4�C  4�  5�J  5�  6 ()%  K�  �  �     )GT  P�  A  �    �  *@  �  �  +h  �  +#  �   �  ,a  p!   ��  �  -h  �  �  �  .�  �� �!   �	  +	  /�  � 0�!1� �   .�  /� �!!   �F	  {	  /�  � 2�  �!   �q	  3�  �� 4�! 5�!�   6U  =�	   �  6�   >�	  6B  ?�	  6�  E�	   �  6B   F�	  6C  G�	  6e  H�	  68  I�	  6�  J�	  6

  X�	   �  6�  Y�	  6�
  Z�	  7�   `&
  �  6�  f7
   �  6�  g7
  6�  h7
  6�  n`
   �  6�	  o`
  6�  p`
  6H  v�
     6`  w�
  6w  x�
  6   y�
  6~  �
     6   ��
  6�  ��
  6  ��
  6�   ��
  6�  ��
  6�	  ��
  6�  �     6  �  6  �  6�  �  6�  �L   %  6�  �L  6�  �L  6�  �L  6m  ��   0  6	  ��  62	  ��  6�  ��  69  ��  6[  ��   ;  6J  ��  6�  ��  67  ��  6�  ��   F  6I	  ��  6$	  ��  6�   �    Q  6N  �   6p  �=   \  6�  �=  6:  �=  6�  �=  6d   �=  6�  �~   g  6  �~  6�  �~  6�	  ѧ   r  6�  ҧ  6  ��   }  6�  ��  6�  ��  6�  ��  6+  ��   �  6�  ��  6�   ��  6  �"   �  6�
  �"  6�  �"  6  �K   �  6   �K  6F  �K  6�  �t   �  6�  �t  6�  �t  6D  O�   �  6�  P�  61  Q�  6�  W�   �  6^  X�  6�  3�   �  6�  4�  6�   8    �  6�  9   6l	  =  �  6N  >  6^  ?  6L  @  6a  DR  �  6B  ER  6�	  FR  6  GR  6  HR  6y  IR  6�   �     6�  !�  8�  8�  8�  9�  �1  �    �   EK L� � �b xJ     S� �  �  �x (>   �p  H   �  �x b3   std  8  @	  5(	  6U
  7o
  �S L%  0_� �K  0w  1�  2�  3�  51  6G  7]  8s  :�  ;�  <  =  ?�  @�  Be  C�  D�  E�  G<  HR  Ih  J~  L�  M�  N  O&  Q�  R�  	v  6  
x  K  �  M�   x  O�  �  8  �   �  Qw  �  �  8   �  R  �  �  8     T8  �  �  �  >   x  Z�    8   x  \    8  D   x  _,  7  8     x  cG  R  8  J   �  p�  P  j  u  8  D   �  t�  P  �  �  8  J   �  {�  �  8  =   n	 ~%  �  �  8  P   �  ��    �  �  >   �  �h  V    >    j   :j  �  �`  � #  �?  �D  W  3�  �4  �$  q-  c=  o'  �5   �%  � �8  �X)  ��%  ��  �aO  �Y=  � P  �� �C  ��wS  ��O  � �?  ��5  �� 
$ g   )W  �   �U  �A  �8  �P   EH  �� �4  �-  O   �7  (  �Q  G  �� b4 �  �P  �8  �4  P  6  dec P  t-  P  hex P  r'  P  < P   oct P  @� P  �[)  P   �%  "P   �  &P   dO  )P   \=  ,P   �P  /P    �C  3P   @zS  6P  ��O  9P  J�?  <P  �  J   (  Qf  K  �Q  Vf  O  Yf   �9  i�  in w�  �  out z�    *  K8  �  8  8   �   !	[ O�   �   "�p 	?]u �  
	   #!�  
q�  =  $!T  H   $]T  %   �  %   
	  6      =  %int (  �  #  �� &�  �  p  �  �  �  �  �O �  o  �O �  �	  pW   ,   qW  !=    "%     #R  ` &�  ` 'p  �^ (�  �^ )�  �T *=  �T +,   iY ,R  hY -%   �e 0�  �e 1p  [ 2=  [ 3,   Q 4=  Q 5,   �_ 6R  �_ 7%   �] :=  �] ;,   �Q >R  �Q ?%   .  <�  `  D=  �  W�  �  _�  �  e=  t   m=  a  u=    ~=  �  �=  3  �=  �  �=  H  �=  y  �=    �=  s  �=  T   �=  �  �=  F  �=  �  �=  �  �=    �=  V  �=  'H   �  (s  Ne  �  Ve  \	  2=  o  7=  �  <=  �  C=  �  =  '		  )'	  H   *pO qO !	  +�  8U
  �{  �   ]�  �  \�   �  �D  !�  �3  "�  U>  #�  &�  $�  �  %�  �*  &�   ڡ  'H   $�U  (H   %TL  )H   &�I  *H   'Q  +H   (�C  ,H   )�J  -H   *1  .�  ,o(  /H   0�U  0H   1PL  1H   2�I  2H   3Q  3H   4�C  4H   5�J  5H   6  )%  K�  o
  =  
	   ,GT  Pz
  '(	  	$   '  �  $,�   --  "�� 1�� �
  
	  
	   -V� Hp� =  �
  �  �   �    .A� ez =  �  �   
	  O     �� �� �  	2*  7*  /8�    Ye �[ 'j  '  0  1j  0j  '(    
	  2�  �  3__a K8  3__b K8   4�
  �!~   �  5��  1
	  � 5{�  1
	  �6 J 7R'  4�  �� 8�*  6  ��~9�� 8�  k:__e :  S;+"�  ;>"�    <H     =�  k   �  4�
  @"g   ��  5��  H�  � 5f� H�   �5\;  H�   �6 J 8� M%   ��,�%�9��  R=  7��  S�  �� 7R'  T�   (� ;l"�  ;�"�    4�
  �"  �~  5��  e�  � 5f� e�   �5-  e
	  �>�| fO   Q� 6@J ?__d h�  �� ?__s i
	  �� 7_X jc  �� @`J M  ?__v x
	  *�  A|#4   s  7R'  �8  =� ;�#"   ;�#�    9U  =�   �  9�   >�  9B  ?�  9�  E�   �  9B   F�  9C  G�  9e  H�  98  I�  9�  J�  9

  X    �  9�  Y   9�
  Z   B�   `)  �  9�  f:   �  9�  g:  9�  h:  9�  nc   �  9�	  oc  9�  pc  9H  v�   �  9`  w�  9w  x�  9   y�  9~  �     9   ��  9�  ��  9  ��  9�   ��  9�  ��  9�	  ��  9�  �     9  �  9  �  9�  �  9�  �O     9�  �O  9�  �O  9�  �O  9m  ��   #  9	  ��  92	  ��  9�  ��  99  ��  9[  ��   .  9J  ��  9�  ��  97  ��  9�  ��   9  9I	  ��  9$	  ��  9�   �#   D  9N  �#  9p  �@   O  9�  �@  9:  �@  9�  �@  9d   �@  9�  Ɂ   Z  9  ʁ  9�  ˁ  9�	  Ѫ   e  9�  Ҫ  9  ��   p  9�  ��  9�  ��  9�  ��  9+  ��   {  9�  ��  9�   ��  9  �%   �  9�
  �%  9�  �%  9  �N   �  9   �N  9F  �N  9�  �w   �  9�  �w  9�  �w  9D  O�   �  9�  P�  91  Q�  9�  W�   �  9^  X�  9�  3�   �  9�  4�  9�   8   �  9�  9  9l	  =   �  9N  >   9^  ?   9L  @   9a  DU  �  9B  EU  9�	  FU  9  GU  9  HU  9y  IU  9�   �   �  9�  !�  C�  D�d  �  �  	  �    �C   O >� d� �b (L     g std * R$  v  6�  x  K�  �  MR$   x  Ob   m   T$  R$   	�  Qw  �   �   T$   	�  R  �   �   T$   
  T8  R$  �   �   Z$   x  Z�   �   T$   x  \�   �   T$  `$   x  _�     T$  �   x  c  #  T$  k$   �  p�  q$  ;  F  T$  `$   �  t�  q$  ^  i  T$  k$   �  {y  �  T$  w$   n	 ~%  �  �  T$  q$   �  ��  ~$  �  �  Z$   �  �h  �$  �  Z$    ;    :;   �  	�f$  � �  G�  c�S L%  0@�+  �=  
��  �b  
��(  Fe  
�w$  �3  
�=  X  �+  �+   (  eq 
�<-  ~$  z  �+  �+   lt 
��1  ~$  �  �+  �+   ��  
eF  w$  �  �+  �+  �   �K  
�9  �  �  �+   �(  

!  �+  �  �+  �  �+   1  
�A  �+    �+  �+  �   �5  
�'  �+  A  �+  �+  �   �3  
�A  �+  e  �+  �  (   +  
:  (    �+   3  �C  
 �P  3  �  �+   �B  
$6  ~$  �  �+  �+   eof 
(�:  3  ?  
,N0  3  �+    _� 	��$  0)  1")  28)  3N)  5�)  6�)  7�)  8�)  :Y)  ;o)  <�)  =�)  ?*  @	*  B)  C)  D-)  EC)  G�)  H�)  I�)  J�)  Ld)  Mz)  N�)  O�)  Q**  R*  �?  	��$  K  \>  �$   �e  _�  �4  c�+  �J  d�+  ��  q    �+   ��  s  &  �+  �+   W  y2  �+  w$    �  5,  60-  7J-  �J  p�  �B  �   �   !%  '+   "�B  �  �  k-  '+  �+   #�B  �  k-  w$    �e  y�  $[V  �  �  !�G  !d   <  x�  �4  {�  �J  |�  �J  =&  `S  �\(  ~J  ��  �J  ��  �%  �i  �K  ��   I  ��  :!  �[-   %H  �   8   %�3  2�  %�G  7�+  %t3  B�-  &�'  ��O  �-  
V  ��N  ~$  �  �  �-   
3  �o+  ~$  �  �  �-   	�P  ��O  �  �  }-   	�M  ��P      }-   	�,  �-  *  5  }-  �   
�+  ��R  '+  L  R  }-   
3  �   '+  i  y  }-  �+  �+   �/  !�B  }-  �  �  �  �+   	�O  �|6  �  �  }-  �+   '(  ��6  �  �  }-  �+   (�   �-  '+  �  �  }-   )�1  o�*  '+    }-  �+  �    (�A  $n%  '+  5  ;  q-   (�A  (�I  '+  S  ^  w-  '+   ("A  ,�%  }-  v  |  q-   (�1  2E)    �  �  q-   (�/  6;&    �  �  q-   '�>  :�>  �  �  w-   (S  A:2  �  �  �  q-  �  �+   '�#  K�(  	  #	  q-  �  �  �+   (9  S>$  �  ;	  K	  q-  �  �   (-U  [�7  ~$  c	  n	  q-  �+   *�5  d�-  �	  '+  �+  �   *	1  m�P  �	  '+  �+  �   *�3  v\-  �	  '+  �  �(   *nU  ��-  �	  '+       *nU  �nG  
  '+       *nU  ��   .
  '+  '+  '+   *nU  �IP  N
  '+  �+  �+   �J  �rR  w$  m
  �  �   '�=  ��H  �
  �
  w-  �  �  �   'V  �)  �
  �
  w-   +�'  �D*  �-  ,�0  ��
  �
  w-   -�0  ��
  �
  w-  �+   ,�0  �    w-  �-   ,�0  �   5  w-  �-  �  �   ,�0  �F  `  w-  �-  �  �  �+   ,�0  �q  �  w-  �+  �  �+   ,�0  ��  �  w-  �+  �+   ,�0  ��  �  w-  �  �(  �+   ,�0   �  �  w-  �-   ,�0  �  
  w-  �  �+   ,�0  "  &  w-  w$   .�  *,Q  �-  ?  J  w-  �-   .�  2�G  �-  c  n  w-  �+   .�  =�%  �-  �  �  w-  �(   .�  Mo_ �-  �  �  w-  �-   .�  Y.c �-  �  �  w-  �   .S� f�&    �  �  w-   .S� q�>        q-   /end y<    1  7  w-   /end �6;    P  V  q-   .I ��$  ,  o  u  w-   .I ��7     �  �  q-   .��  �lC  ,  �  �  w-   .��  �CM     �  �  q-   .)^ �^\   �  �  q-   .%] ��a   
    q-   .hf �*]    )  /  q-   .wY �Je    H  N  q-   .r ��R  �  g  m  q-   .�K  �r5  �  �  �  q-   .�3  �j=  �  �  �  q-   0�� ��  �  �  w-  �  �(   0�� ��F  �  �  w-  �   0be  VT     w-   .I  v  �  $  *  q-   0�E  &|U  ?  J  w-  �   0�1  -�  _  e  w-   .�� 5�?  ~$  ~  �  q-   .�:  D�6  �  �  �  q-  �   .�:  UW  �  �  �  w-  �   /at k
/  �  �  �  q-  �   /at ��7  �      w-  �   .��  ��O �  +  1  w-   .��  �}Y �  J  P  q-   .�G  �@\ �  i  o  w-   .�G  �e �  �  �  q-   .�F  ��/  �-  �  �  w-  �-   .�F  �k:  �-  �  �  w-  �+   .�F  ��H  �-  �  �  w-  �(   .�F  �x` �-      w-  �   .@  �A:  �-  7  B  w-  �-   .@  ��1  �-  [  p  w-  �-  �  �   .@  ��D  �-  �  �  w-  �+  �   .@  ��*  �-  �  �  w-  �+   .@  �6  �-  �  �  w-  �  �(   .@  �] �-  �  
  w-  �   0�G  -aN    *  w-  �(   .�3  <b*  �-  C  N  w-  �-   .�3  Ipf �-  g  r  w-  �-   .�3  ^ 2  �-  �  �  w-  �-  �  �   .�3  n�=  �-  �  �  w-  �+  �   .�3  z�T  �-  �  �  w-  �+   .�3  � @  �-      w-  �  �(   .�3  ��a �-  /  :  w-  �   0� ��E  O  d  w-    �  �(   0� ��V y  �  w-    �   .� �\+  �-  �  �  w-  �  �-   .� �u>  �-  �  �  w-  �  �-  �  �   .� |=  �-  �    w-  �  �+  �   .� "�@  �-  ,  <  w-  �  �+   .� 9k<  �-  U  j  w-  �  �  �(   .� K�'    �  �  w-    �(   .bL  d�R  �-  �  �  w-  �  �   .bL  t�2    �  �  w-     .bL  �L&    �  	  w-       0H�  �M\   $  w-   .�%  �9F  �-  =  R  w-  �  �  �-   .�%  �|<  �-  k  �  w-  �  �  �-  �  �   .�%  ��T  �-  �  �  w-  �  �  �+  �   .�%  ��A  �-  �  �  w-  �  �  �+   .�%  b>  �-      w-  �  �  �  �(   .�%  3%  �-  7  L  w-      �-   .�%  'V7  �-  e    w-      �+  �   .�%  <�+  �-  �  �  w-      �+   .�%  Q'S  �-  �  �  w-      �  �(   .�%  vj.  �-  �    w-      '+  '+   .�%  ��9  �-  ,  F  w-      �+  �+   .�%  �C  �-  _  y  w-           .�%  �>/  �-  �  �  w-           .�%  �b �-  �  �  w-      �   (�?  ��&  �-  �    w-  �  �  �  �(   (�1  �O  �-  $  >  w-  �  �  �+  �   ,)  �z-  '+  b  �  �(  �+   +E  �3J  '+  �  �  �(  �+   .�5  �)  �  �  �  q-  '+  �  �   0n	 @D  �  �  w-  �-   .W�  �6  �+  �  �  q-   .�A  %�A  �+      q-   .��  ,Z5  �  +  1  q-   .�(  <;  �  J  _  q-  �+  �  �   .�(  I�%  �  x  �  q-  �-  �   .�(  X�5  �  �  �  q-  �+  �   .�(  i^   �  �  �  q-  �(  �   .�(  v�S  �  �    q-  �-  �   .�(  �K  �    1  q-  �+  �  �   .�(  �o?  �  J  Z  q-  �+  �   .�(  �J5  �  s  �  q-  �(  �   .NW  ��Q  �  �  �  q-  �-  �   .NW  ��I  �  �  �  q-  �+  �  �   .NW  ��,  �  �    q-  �+  �   .NW  ��;  �    ,  q-  �(  �   .�S  ��I  �  E  U  q-  �-  �   .�S  T?  �  n  �  q-  �+  �  �   .�S  05  �  �  �  q-  �+  �   .�S  $S:  �  �  �  q-  �(  �   .�>  2hL  �  �  �  q-  �-  �   .�>  CUB  �    ,  q-  �+  �  �   .�>  Q�2  �  E  U  q-  �+  �   .�>  b�K  �  n  ~  q-  �(  �   .�4  qT  �  �  �  q-  �-  �   .�4  ��K  �  �  �  q-  �+  �  �   .�4  ��5  �  �  �  q-  �+  �   .�4  �N.  �    '  q-  �(  �   .U+  �)  X  @  P  q-  �  �   .��  �!1  w$  i  t  q-  �-   .��  ��T  w$  �  �  q-  �  �  �-   .��  ��O  w$  �  �  q-  �  �  �-  �  �   .��  	;.  w$  �  �  q-  �+   .��  (	�B  w$    ,  q-  �  �  �+   .��  C	�,  w$  E  _  q-  �  �  �+  �   i  1!T  �(  2�E    2�F  �   � >X  �&  �7  X  Qf /z  �J  6�+  t :�   �e  5�  �x ;�  `S  7�+  3�w >�    S/  �  �   �w B    S/   r G�i �  /  5  Y/   S� K�m �  M  S  Y/   4end O;u �  k  q  Y/   5_E �(   � '6��  )<�-  =�-  >�-  @R.  A].  Bw.  C�.  D�.  E�.  F�.  G/  H/  Gz <�  7_V2 �8��       Y� �x w)!  9~ �w$   9z �;/  3�x y:   @   A/   3�x |O   _   A/  w$  G/   	�3  �Nz r   �   A/  w$  G/   	�1  ��y �   �   A/   
~ ��� w$  �   �   M/   
�| ��| G/  �   �   M/   
} ��y .!  �   �   M/   
9� ��y �  	!  !  M/   :�  �� ~$  "!  M/       �� �;"  ~ �w$   z �;/  �� �b!  h!  _/   �� �x!  �!  _/  w$  G/   �3  ҁ{ �!  �!  _/  w$  G/   �1  ��} �!  �!  _/   ~ ��{ w$  �!  �!  e/   �| �} G/  �!  "  e/   9� ��x �  "   "  e/   ;�  �y ~$  4"  e/    �  .!  6yy a6o� d6� hPa(  Q�(  Ra(  Sa(  Ta(  <�� 8�"  =#�  =� =�� =�� =�� =)�  >�~ @�"  =�| =�y =�~ =  ד  �#  ��  ��  � �'+  �4  ��+  1{�  '+   ?N| ^�#  �#  �#   )� `   @N| cC#  N#  e0      A8� K#  c#  n#  e0  w$   B(� N�� �+  #  �#  �#  k0   ,� m�� k/  �#  k0    �p #  �� &1 H�{ G/  C%�  e �  �#  �  D	[ O�#     D6y ) $   z  EIc  1$   �  E& j&$   E"  E�~ k9$   N"  E{ lL$   W"   FG;   G�  H�  I�  J;   H;   Kint L�  G�  L�  L�  Lo  L�  L�  L�  L�	  L(  L#  $   ��(  �  $,�  -�  K  :8&  �e  =�  � ?'+  "  @�+  �4  A�+  �J  B�+  �A  OB%  H%  �+   �A  QX%  c%  �+  �+   �A  Vs%  ~%  �+  w$   �
 Y51  %  �%  �%  �+  %   �
 ]�R  %  �%  �%  �+  &%   � c?  %  �%  �%  �+  �$  �+   _ m.    &  &  �+  %  �$   �3  q89  �$  (&  .&  �+   5_Tp �(   �$  MZD  �\(  NF�  �'+   O��  ��"  O�4  ��"  O� ��"  ,��  ��&  �&  H0   -��  ��&  �&  H0  N0   .*  ��}  e&  �&  �&  Y0   .Ư  �?s  r&  �&  �&  Y0   .�F  �Ϭ  _0  	'  '  H0   .�F  ��  =&  ('  3'  H0  w$   .a�  �
�  _0  L'  R'  H0   .a�   ��  =&  k'  v'  H0  w$   .�:  ,�  e&  �'  �'  Y0  X&   .�F  		n  _0  �'  �'  H0  X&   .(*  ��  =&  �'  �'  Y0  X&   . I  h�  _0  �'  (  H0  X&   .�O  7k  =&  (  *(  Y0  X&   .WC  ]�  N0  C(  I(  Y0   1{�  '+  1�  X   8E  <*; 1�(  =�8  =�; =N;  P�= 5�(   a(  =&  QU  A[-  �(  �0  w$   R9+  N[-  �0  w$    L�� L�� L�� 2*  7�(  S8   _�  ԋ$  L�  �  !�$  �  !�$  �O !�$  �O !�$  pW  ! �$  qW  !!w$    !"�$    !#�$  ` !&�$  ` !'�$  �^ !(�$  �^ !)�$  �T !*w$  �T !+�$  iY !,�$  hY !-�$  �e !0�$  �e !1�$  [ !2w$  [ !3�$  Q !4w$  Q !5�$  �_ !6�$  �_ !7�$  �] !:w$  �] !;�$  �Q !>�$  �Q !?�$  .  "<8)  `  "Dw$  �  "W8)  �  "_C)  �  "ew$  t   "mw$  a  "uw$    "~w$  �  "�w$  3  "�w$  �  "�w$  H  "�w$  y  "�w$    "�w$  s  "�w$  T   "�w$  �  "�w$  F  "�w$  �  "�w$  �  "�w$    "�w$  V  "�w$  G�(  L�  s  #N)  �  #V)  \	  $2w$  o  $7w$  �  $<w$  �  $Cw$  �  %w$  G�+  TG�+  �(  U&pO qO &!�+  H(  HX  GX  G(  H  LYe L�[ H�(  H�+  G�$  H8&  G8&  G�  H>  L  �  8'0-  �{  ''+   ]�  ''+  \�  ' '+  �D  '!'+  �3  '"'+  U>  '#'+  &�  '$'+  �  '%'+  �*  '&'+   ڡ  ''�(  $�U  '(�(  %TL  ')�(  &�I  '*�(  'Q  '+�(  (�C  ',�(  )�J  '-�(  *1  '.'+  ,o(  '/�(  0�U  '0�(  1PL  '1�(  2�I  '2�(  3Q  '3�(  4�C  '4�(  5�J  '5�(  6 V)%  'K'+  J-  w$  �+   WGT  'PU-  G,  �  ( w$  w$  Gd  G�  GX  Gi  Hi  H�  JX  HX  X�$  �-  Y G_  �l  )�$  j�  )#�$  Ztm ,),R.  ,g  ).w$   �  )/w$  �  )0w$  ��  )1w$  ��  )2w$  ��  )3w$  ��  )4w$  �  )5w$  d�  )6w$   ��  )7�$  $~�  )8�+  ( W\�  )>�-  Vѯ  )H�(  w.  �-  �-   V��  )M�-  �.  �.   G�-  V�  )C�-  �.  �.   G�-  V#�  )a'+  �.  �.   G�.  �-  V�� )f'+  �.  �.   G�.  �-  V��  )W�.  /  �.   V[v  )\�.  /  �.   V��  )R�(  ;/  '+  �(  �+  �.   G�  G   H�  G)!  G�  G;"  G.!  G@"  H)!  [A0  \�     00        ]� �/  �/  q0  w0   ]� �/  �/  q0  }0   ]� �/  �/  q0   ^H�   �+  v/  �/  �/  �0   ^9� #�  v/  0  0  �0  w$   _� v/  $0  q0  w$    v/  `�� =}0   Sq/  G=&  HT0  '+  G�(  H=&  G#  G�#  Gv/  Jv/  H00  G00  G[-  a�(  �0  bXF  A�0  b\;  Aw$  cd�T  C[-    e  �0  �0  fh  �0   q-  a�  �0  cg__p �R$    h0  1  1  fh  1  f#  f-   q0  a�(  ;1  bXF  N�0  b\;  Nw$   e�  I1  ^1  fh  ^1  i__a �c1   }-  �+  eN#  v1  �1  fh  �1  f#  f-   e0  a�  �1  j__s 
�+   e�   �1  �1  fh  �1   M/  e�   �1  �1  fh  �1   e2%  �1  �1  fh  �1   �+  e�  2  2  fh  2   �+  ec%  "2  52  fh  �1  f#  f-   e&  C2  V2  fh  2  f#  f-   eH%  d2  s2  fh  �1  s2   �+  e  �2  �2  fh  2  i__a s�2   �+  e  �2  �2  fh  �0   e^  �2  �2  fh  �0   k�  �2  �2  fh  �2  f#  f-   k-  e�   3  3  fh  �1   e�  3  )3  fh  �0   e
  73  J3  fh  J3  f#  f-   w-  e�  ]3  3  fh  �2  lv�  '+  j__a 3   �+  m�
  e5  �3  �3  fh  ^1   e�
  �3  �3  fh  J3   eJ  �3  �3  fh  J3  j__s 2�+   n�/  �#   ��3  4  oh  4  �  �0  p�0  �#   �4  54  q1  � r�#s� �   p�0  �#!   �L4  �4  q1  � t�0  �#   v4  u1  P� v�# w$C   xh1  L� $   ��4  �4  qv1  � r$s� �   xh1  ��  $!   ��4  5  qv1  � th1  ($   K�4  uv1  o� v4$ wA$C   e�/  5  85  fh  4  b�} #w$  cd��  %�  cy73     e�  F5  \5  fh  J3  j__s z�+   zn#  P$o  �s5  �9  oh  �9  � {�2  b$�J N�8  u3  �� |5  s$�J �u5  �� u5  m� }�J ~$5  t�3  v$   %6  u�3  �� O3  v$   �yr3  uf3  �� u]3  ��   t�3  �$   )^6  u�3  6� u�3  N� 85  �$   3uO5  6� uF5  N� ��$�    t�3  �$   ,�6  u�3  {� u�3  �� 85  �$   3uO5  {� uF5  �� ��$�    {�3  �$�J 57  u�3  �� u�3  �� �85  �$�J 3uO5  �� uF5  �� �C%�    t�3  P%    2X7  u�3  � u�3  � 85  P%    3uO5  � uF5  � �c%�    t�3  p%   /�7  u�3  J� u�3  b� 85  p%   3uO5  J� uF5  b� ��%�    ��%7   q73  ud���2  �%   #�7  q�2  ud��0  �%   -q�0  ud�  ;1  �%/   #qR1  uc�uI1  �� ��%   uR1  �� uI1  �� {1  �% K ��8  �/1  u$1  �� |�0  �% K V��0  u�0  �� } K ��0  S   ��%�        {3  �$K N�8  u3  � ��0  �$K u�0  �   {)3  �$0K N�9  u73  � ��2  �$HK #
9  u�2  �  �;1  �$`K #uR1  "� uI1  D� ��$'   uR1  b� uI1  �� {1  �$xK ��9  u/1  �� u$1  �� |�0  �$xK Vu�0  �� u�0  �� }xK ��0  ��    ��$�     ��%"C   k0  p5  �%  ��9  �<  q5  �q5  ���K �<  �$5  � t�3  �%   %>:  u�3  �� O3  �%   �yr3  uf3  �� u]3  ��   t�3  �%   )�:  u�3  �� u�3  �� 85  �%   3uO5  �� uF5  �� ��%�    {�3  �%�K 5�:  u�3   � u�3  � �85  �%�K 3uO5   � uF5  � �p&�    t�3  &   28;  u�3  8� u�3  P� 85  &   3uO5  8� uF5  P� � &�    t�3  5&   ,�;  u�3  p� u�3  �� 85  5&   3uO5  p� uF5  �� �E&�    t�3  �&   /�;  u�3  �� u�3  �� 85  �&   3uO5  �� uF5  �� ��&�    ��&6   u73  �� ��2  �&   #*<  u�2  �� �0  �&   -u�0  ��   ;1  �&/   #qR1  ug�uI1   � ��&   uR1  � uI1  K� {1  �&�K ��<  �/1  u$1  ^� |�0  �&�K V��0  u�0  ^� }�K ��0  S   ��&�      ��&"C   a50  �<  cdF� ?00    ��#  �&T   �@=  |�<  �&L I}L ��<  �D��&6C  �'PC  �('`C     �U  "=M=   5*  ��   ">M=  �B  "?M=  ��  "Ey=   @*  �B   "Fy=  �C  "Gy=  �e  "Hy=  �8  "Iy=  ��  "Jy=  �

  "X�=   K*  ��  "Y�=  ��
  "Z�=  ��   "`�=  V*  ��  "f
>   a*  ��  "g
>  ��  "h
>  ��  "n6>   l*  ��	  "o6>  ��  "p6>  �H  "vb>   w*  �`  "wb>  �w  "xb>  �   "yb>  �~  "�>   �*  �   "��>  ��  "��>  �  "��>  ��   "��>  ��  "��>  ��	  "��>  ��  "��>   �*  �  "��>  �  "��>  ��  "��>  ��  "�4?   �*  ��  "�4?  ��  "�4?  ��  "�4?  �m  "�m?   �*  �	  "�m?  �2	  "�m?  ��  "�m?  �9  "�m?  �[  "��?   �*  �J  "��?  ��  "��?  �7  "��?  ��  "��?   �*  �I	  "��?  �$	  "��?  ��   "�@   �*  �N  "�@  �p  "�7@   �*  ��  "�7@  �:  "�7@  ��  "�7@  �d   "�7@  ��  "�}@   �*  �  "�}@  ��  "�}@  ��	  "ѩ@   �*  ��  "ҩ@  �  "��@   �*  ��  "��@  ��  "��@  ��  "��@  �+  "�A   �*  ��  "�A  ��   "�A  �  "�-A   +  ��
  "�-A  ��  "�-A  �  "�YA   +  �   "�YA  �F  "�YA  ��  "�A   +  ��  "�A  ��  "��A  �D  #O�A   4+  ��  #P�A  �1  #Q�A  ��  #W�A   ?+  �^  #X�A  ��  $3�A   J+  ��  $4�A  ��   $8B   U+  ��  $9B  �l	  $=:B  `+  �N  $>:B  �^  $?:B  �L  $@:B  �a  $DsB  k+  �B  $EsB  ��	  $FsB  �  $GsB  �  $HsB  �y  $IsB  ��  % �B   v+  ��  %!�B  ��� R$  ��(   ��#  ��#  �$  �$  �+$  �>$  �  �1  "C  R$   �>  Y  6C  R$   �e= w$  JC  JC   G�$  �Y< `C  JC   �� w$  ~C  ~C  R$  R$   G�C  �R$     =   �W �� �� �b �L     � (  _� �7   �  #  �� �  std   5%  R5%  Uh%  [�%  \�%  @q(  v  61  x  K+  	�  M(   
x  O�   �   |(  (   �  Qw  �   �   |(   �  R  �   �   |(     T8  (      �(   x  Z  !  |(   x  \1  <  |(  �(   x  _L  W  |(  8   x  cg  r  |(  �(   �  p�  �(  �  �  |(  �(   �  t�  �(  �  �  |(  �(   �  {�  �  |(  O%   n	 ~%  �  �  |(  �(   �  ��  �(  
    �(   �  �h  �(  $  �(    �    :�   �  �L   � C  �S !L%  0�=  �$  �b  �a%  Fe  �O%  �3  �=  �  e,  k,   h  eq �<-  �(  �  k,  k,   lt ��1  �(  �  k,  k,   ��  eF  O%  �  q,  q,  $   �K  �9  $    q,   �(  
!  q,  9  q,  $  k,   1  �A  w,  ]  w,  q,  $   �5  �'  w,  �  w,  q,  $   �3  �A  w,  �  w,  $  h   +  :  h  �  },   s  �C   �P  s  �  k,   �B  $6  �(  �  },  },   eof (�:  s  ?  ,N0  s  },    _� �7   	0�%  	1�%  	2&  	33&  	5�&  	6�&  	7�&  	8�&  	:>&  	;T&  	<j&  	=�&  	?'  	@�&  	B�%  	C�%  	D&  	E!&  	G�&  	H�&  	I�&  	J�&  	LI&  	M_&  	Nu&  	O�&  	Q'  	R�&  �?  �%   K  
\~  �(   �e  
_$  �4  
c�,  �J  
d�,  ��  
qE  K  �,   ��  
s[  f  �,  �,    W  
yr  �,  O%    �  5�,  6�-  7	.  �J  p�  !�B  �  "�   #%  }%   $�B  �  0.  }%  �,    �e  y  %[V  �  �  #�G  !�   <  x�  �4  {  �J  |)  �J  *  `S  �9,  ~J  ��  �J  ��  �%  ��  	�K  ��   	I  ��  	:!  �.   %H  �E  "`   &�3  2�  &�G  7\%  &t3  B`.  '�'  ��O  H.  V  ��N  �(  �  �  k.   3  �o+  �(      k.   �P  ��O     &  B.   �M  ��P  9  ?  B.   �,  �-  R  ]  B.  �   �+  ��R  }%  t  z  B.   3  �   }%  �  �  B.  �,  �,   �/  !�B  B.  �  �  �  �,   �O  �|6  �  �  B.  �,   ((  ��6  �    B.  �,   )�   �-  }%       B.   *�1  o�*  }%  4  B.  �,  �    )�A  $n%  }%  ]  c  6.   )�A  (�I  }%  {  �  <.  }%   )"A  ,�%  B.  �  �  6.   )�1  2E)  0  �  �  6.   )�/  6;&  0  �  �  6.   (�>  :�>  �  �  <.   )S  A:2  �  	  "	  6.  �  V%   (�#  K�(  6	  K	  6.  �  �  V%   )9  S>$  �  c	  s	  6.  �  �   )-U  [�7  �(  �	  �	  6.  V%   +�5  d�-  �	  }%  V%  �   +	1  m�P  �	  }%  V%  �   +�3  v\-  �	  }%  �  a%   +nU  ��-  
  }%  0  0   +nU  �nG  6
  }%  <  <   +nU  ��   V
  }%  }%  }%   +nU  �IP  v
  }%  V%  V%   �J  �rR  O%  �
  �  �   (�=  ��H  �
  �
  <.  �  �  �   (V  �)  �
  �
  <.   ,�'  �D*  H.  -�0  ��
  �
  <.   .�0  �    <.  �,   -�0  �,  7  <.  N.   -�0  �H  ]  <.  N.  �  �   -�0  �n  �  <.  N.  �  �  �,   -�0  ��  �  <.  V%  �  �,   -�0  ��  �  <.  V%  �,   -�0  ��  �  <.  �  a%  �,   -�0       <.  T.   -�0  "  2  <.  �  �,   -�0  "C  N  <.  O%   /�  *,Q  Z.  g  r  <.  N.   /�  2�G  Z.  �  �  <.  V%   /�  =�%  Z.  �  �  <.  a%   /�  Mo_ Z.  �  �  <.  T.   /�  Y.c Z.  �    <.  �   /S� f�&  0    !  <.   /S� q�>  <  :  @  6.   0end y<  0  Y  _  <.   0end �6;  <  x  ~  6.   /I ��$  T  �  �  <.   /I ��7  H  �  �  6.   /��  �lC  T  �  �  <.   /��  �CM  H  �  �  6.   /)^ �^\ <      6.   /%] ��a <  2  8  6.   /hf �*] H  Q  W  6.   /wY �Je H  p  v  6.   /r ��R  �  �  �  6.   /�K  �r5  �  �  �  6.   /�3  �j=  �  �  �  6.   1�� ��  �  �  <.  �  a%   1�� ��F      <.  �   1be  VT -  3  <.   /I  v  �  L  R  6.   1�E  &|U  g  r  <.  �   1�1  -�  �  �  <.   /�� 5�?  �(  �  �  6.   /�:  D�6  $  �  �  6.  �   /�:  UW    �  �  <.  �   0at k
/  $      6.  �   0at ��7    /  :  <.  �   /��  ��O   S  Y  <.   /��  �}Y $  r  x  6.   /�G  �@\   �  �  <.   /�G  �e $  �  �  6.   /�F  ��/  Z.  �  �  <.  N.   /�F  �k:  Z.  �  �  <.  V%   /�F  ��H  Z.    "  <.  a%   /�F  �x` Z.  ;  F  <.  �   /@  �A:  Z.  _  j  <.  N.   /@  ��1  Z.  �  �  <.  N.  �  �   /@  ��D  Z.  �  �  <.  V%  �   /@  ��*  Z.  �  �  <.  V%   /@  �6  Z.  �    <.  �  a%   /@  �] Z.  '  2  <.  �   1�G  -aN  G  R  <.  a%   /�3  <b*  Z.  k  v  <.  N.   /�3  Ipf Z.  �  �  <.  T.   /�3  ^ 2  Z.  �  �  <.  N.  �  �   /�3  n�=  Z.  �  �  <.  V%  �   /�3  z�T  Z.  
    <.  V%   /�3  � @  Z.  .  >  <.  �  a%   /�3  ��a Z.  W  b  <.  �   1� ��E  w  �  <.  0  �  a%   1� ��V �  �  <.  0  �   /� �\+  Z.  �  �  <.  �  N.   /� �u>  Z.  �    <.  �  N.  �  �   /� |=  Z.  &  ;  <.  �  V%  �   /� "�@  Z.  T  d  <.  �  V%   /� 9k<  Z.  }  �  <.  �  �  a%   /� K�'  0  �  �  <.  0  a%   /bL  d�R  Z.  �  �  <.  �  �   /bL  t�2  0  �    <.  0   /bL  �L&  0  !  1  <.  0  0   1H�  �M\ F  L  <.   /�%  �9F  Z.  e  z  <.  �  �  N.   /�%  �|<  Z.  �  �  <.  �  �  N.  �  �   /�%  ��T  Z.  �  �  <.  �  �  V%  �   /�%  ��A  Z.  �    <.  �  �  V%   /�%  b>  Z.  ,  F  <.  �  �  �  a%   /�%  3%  Z.  _  t  <.  0  0  N.   /�%  'V7  Z.  �  �  <.  0  0  V%  �   /�%  <�+  Z.  �  �  <.  0  0  V%   /�%  Q'S  Z.  �    <.  0  0  �  a%   /�%  vj.  Z.  !  ;  <.  0  0  }%  }%   /�%  ��9  Z.  T  n  <.  0  0  V%  V%   /�%  �C  Z.  �  �  <.  0  0  0  0   /�%  �>/  Z.  �  �  <.  0  0  <  <   /�%  �b Z.  �    <.  0  0  �   )�?  ��&  Z.    4  <.  �  �  �  a%   )�1  �O  Z.  L  f  <.  �  �  V%  �   ,)  �z-  }%  �  �  a%  �,   +E  �3J  }%  �  �  a%  �,   /�5  �)  �  �  �  6.  }%  �  �   1n	 @D  �  �  <.  Z.   /W�  �6  V%      6.   /�A  %�A  V%  4  :  6.   /��  ,Z5    S  Y  6.   /�(  <;  �  r  �  6.  V%  �  �   /�(  I�%  �  �  �  6.  N.  �   /�(  X�5  �  �  �  6.  V%  �   /�(  i^   �  �    6.  a%  �   /�(  v�S  �    +  6.  N.  �   /�(  �K  �  D  Y  6.  V%  �  �   /�(  �o?  �  r  �  6.  V%  �   /�(  �J5  �  �  �  6.  a%  �   /NW  ��Q  �  �  �  6.  N.  �   /NW  ��I  �  �    6.  V%  �  �   /NW  ��,  �    +  6.  V%  �   /NW  ��;  �  D  T  6.  a%  �   /�S  ��I  �  m  }  6.  N.  �   /�S  T?  �  �  �  6.  V%  �  �   /�S  05  �  �  �  6.  V%  �   /�S  $S:  �  �  �  6.  a%  �   /�>  2hL  �    &  6.  N.  �   /�>  CUB  �  ?  T  6.  V%  �  �   /�>  Q�2  �  m  }  6.  V%  �   /�>  b�K  �  �  �  6.  a%  �   /�4  qT  �  �  �  6.  N.  �   /�4  ��K  �  �  �  6.  V%  �  �   /�4  ��5  �    &  6.  V%  �   /�4  �N.  �  ?  O  6.  a%  �   /U+  �)  �  h  x  6.  �  �   /��  �!1  O%  �  �  6.  N.   /��  ��T  O%  �  �  6.  �  �  N.   /��  ��O  O%  �    6.  �  �  N.  �  �   /��  	;.  O%    &  6.  V%   /��  (	�B  O%  ?  T  6.  �  �  V%   /��  C	�,  O%  m  �  6.  �  �  V%  �   �  2!T  a%  3�E  \  3�F  �   �  � >�  �&  �7  �  Qf /�  �J  6V%  	t :�   �e  5$  	�x ;�  `S  7V%  4�w >  .  �.    �   �w B>  D  �.   r G�i �  \  b  �.   S� K�m   z  �  �.   5end O;u   �  �  �.   6_E a%   �  7Y� B�  }!  8S� �0   Y� H�  �  �0   9$� B�  �  �  �0  O%   Y� M      �0  �.   �  N�� �0  0   ;   �0  �.   :H�  Q�� V%  �  [   a   q.   :9� T�� �  �  �   �   q.  O%   :} T=� �"  �  �   �   q.  O%   :v� Xh� �(  �  �   �   q.  O%  �0   :v� ]�� �(  �  !  !  q.  �.  O%   }� `�� �(  /!  :!  q.  �.   U  d�� �(  R!  ]!  q.  �.   2  h� �(  q!  q.  �.    �x w�"  ;~ �O%   ;z �q.  4�x y�!  �!  |.   4�x |�!  �!  |.  O%  �.   �3  �Nz �!  �!  |.  O%  �.   �1  ��y "  "  |.   ~ ��� O%  *"  0"  �.   �| ��| �.  G"  M"  �.   } ��y �"  d"  j"  �.   9� ��y �  �"  �"  �.   <�  �� �(  �"  �.    }!  �� ĳ#  	~ �O%   	z �q.  �� ��"  �"  �.   �� ��"   #  �.  O%  �.   �3  ҁ{ #  $#  �.  O%  �.   �1  ��} 8#  >#  �.   ~ ��{ O%  V#  \#  �.   �| �} �.  t#  z#  �.   9� ��x �  �#  �#  �.   =�  �y �(  �#  �.    �  �"  ד  ��#  ��  ��  � �}%  �4  ��,  2{�  }%   >| 8�$  �$  �$   #)� ;}!  -| >*$  5$  q0  }!   -| AF$  V$  q0  }!  *.   -| Og$  w$  q0  O%  �.   -| S�$  �$  q0  O%  �.  *.   ?o� 8�#  �$  �$  q0  O%   @,� Z� �.  �$  w0    �8 �#  �� AU  �(  %  �0  �0   '� L�� �.  '�| Oy �.  B	[ !O/%   M   C��  EO%  O%  V%  V%   Dint E\%  a%  �  C��  U}%  }%  O%   Ea%  C��  O}%  �%  }%  V%   C��  F,   �%  }%  V%  ,    �  �%  �  �  �%  �  �O �%  o  �O �%  �	  pW   &  �  qW  !O%    ",&  �    #>   ` &�%  ` '�%  �^ (�%  �^ )�%  �T *O%  �T +&  iY ,>   hY -,&  �e 0�%  �e 1�%  [ 2O%  [ 3&  Q 4O%  Q 5&  �_ 6>   �_ 7,&  �] :O%  �] ;&  �Q >>   �Q ?,&  .  <&  `  DO%  �  W&  �  _!&  �  eO%  t   mO%  a  uO%    ~O%  �  �O%  3  �O%  �  �O%  H  �O%  y  �O%    �O%  s  �O%  T   �O%  �  �O%  F  �O%  �  �O%  �  �O%    �O%  V  �O%  �  Fs  N�%  �  V�%  \	  2O%  o  7O%  �  <O%  �  CO%  �  O%  Eh(  GHpO qO !i(  E�   E+  I+  J�   I�   �  EH  $   �D,  �  $,$  -�  K  :*  �e  =$  � ?}%  "  @V%  �4  A�,  �J  B�,  �A  O)  %)  �,   �A  Q5)  @)  �,  �,   �A  VP)  [)  �,  O%   �
 Y51  �(  s)  ~)  �,  �(   �
 ]�R  �(  �)  �)  �,  )   � c?  �(  �)  �)  �,  �(  b(   _ m.   �)  �)  �,  �(  �(   �3  q89  �(  *  *  �,   6_Tp a%   �(  KZD  �9,  LF�  �}%   M��  ��#  M�4  ��#  M� ��#  -��  �m*  s*  T0   .��  ��*  �*  T0  Z0   /*  ��}  B*  �*  �*  e0   /Ư  �?s  O*  �*  �*  e0   /�F  �Ϭ  k0  �*  �*  T0   /�F  ��  *  +  +  T0  O%   /a�  �
�  k0  )+  /+  T0   /a�   ��  *  H+  S+  T0  O%   /�:  ,�  B*  l+  w+  e0  5*   /�F  		n  k0  �+  �+  T0  5*   /(*  ��  *  �+  �+  e0  5*   / I  h�  k0  �+  �+  T0  5*   /�O  7k  *  �+  ,  e0  5*   /WC  ]�  Z0   ,  &,  e0   2{�  }%  2�  �   8E  *   �� �� 2*  7e,  N8U   Ih  I�  E�  Eh  I�  Ye �[ Ia%  I\%  E�(  I*  E*  E�  I~    �  8�-  	�{  }%   	]�  }%  	\�   }%  	�D  !}%  	�3  "}%  	U>  #}%  	&�  $}%  	�  %}%  	�*  &}%   	ڡ  'a%  $	�U  (a%  %	TL  )a%  &	�I  *a%  '	Q  +a%  (	�C  ,a%  )	�J  -a%  *	1  .}%  ,	o(  /a%  0	�U  0a%  1	PL  1a%  2	�I  2a%  3	Q  3a%  4	�C  4a%  5	�J  5a%  6 C)%  K}%  	.  O%  V%   OGT  P.  E�,  �   O%  O%  I�  E�  E�  E�  E�  I�  I�  J�  I�  P7   k.  Q E�  E�  q.  E}!  I�  E�"  E�  E�#  E�"  E�#  I�"  RM0  !�  S�� 2�  r/  "�   T�� �.  �.  �0  �0   T�� �.  �.  �0  �0   T�� /  /  �0   UH�  5V%  �.  ,/  2/  �0   U9� 9�  �.  M/  X/  �0  O%   V�� �.  f/  �0  O%    �.  S� #�  10  "�   T� �/  �/  �0  �0   T� �/  �/  �0  �0   T� �/  �/  �0   UH�  &V%  w/  �/  �/  �0   U9� *�  w/  0  0  �0  O%   V� w/  %0  �0  O%    w/  W9� A10  W]� Br/   N �.  E*  I`0  }%  E>,  I*  E�#  E�$  XO%  �0  Y E�0  Z�5  }0  E�  I�  I�#  E�.  J�.  Ir/  Er/  Ew/  Jw/  I10  E10  [�$  �0  �0  \h  �0  \#  %.   q0  ["  1  1  \h  1   �.  [0"  +1  51  \h  1   [:!  C1  X1  \h  w.  ]�< dX1   �.  [�"  k1  �1  \h  �1  ^__v �O%  ]=8 ɐ1   �.  �.  [>#  �1  �1  \h  �1   �.  [\#  �1  �1  \h  �1   _�$  �1  `\C  �1  `?)  �1   �0  �0  [�  2  2  \h  2  \#  %.   �0  aX/  2-2  @2  \h  @2  \#  %.   �0  a0  #U2  h2  \h  h2  \#  %.   �0  [)  {2  �2  \h  �2   �,  [5  �2  �2  \h  �2   �,  [@)  �2  �2  \h  �2  \#  %.   [f  �2  �2  \h  �2  \#  %.   b^�  
3  ]w  eO%  ]-�  eO%   c�/  @'   �!3  .3  dh  .3  �  �0  c/  P'   �J3  W3  dh  W3  �  �0  [�   j3  3  \h  w.  ^__i TO%   e\3  =� `'   ��3  �3  fj3  �fs3  �g]1  d'   Uf1  �ft1  �fk1  �   c�   �'*   ��3  4  dh  w.  � h�� ]4  �i__i ]O%  � �.  j2  �'   �/4  84  f-2  �  jE2  �'   �O4  X4  fU2  �  j2  �'   �o4  �4  f-2  � k�'�<  l� �   jE2  �'   ��4  �4  fU2  � k�'�<  l� �   c2/  �')   ��4  �4  dh  W3  �ii 9O%  �m(h%  n( c�/   ()   �5  85  dh  .3  �ii *O%  �m1(h%  n@( e�0  �� P(   �S5  j5  f�0  � o_(l� �   e�0  �� `(!   ��5  �5  f�0  � p�0  h(   8�5  q�0  s� nt( r�(�<   s�   �(Y   ��5  U6  dh  w.  � i__i XO%  �h�� YU6  �t\3  �(   Z66  us3  uj3  g]1  �(   Uu1  ut1  uk1    v�1  �(pL Zq�1  �� u�1    �0  e�1  C� �(   �u6  ~6  f2  �  e�1  ��  )   ��6  �6  f2  � k)�<  l� �   w%  )   �w%   )   �xM"  a0)J   ��6  E7  dh  1  �g\3  N)   bqs3  �� qj3  �� g]1  N)   Uq1  �� qt1  �� qk1  ��    y4� ��2   ��7  g�2  ��+   ez�2  {�2  ��mǁ�<  mށ�<    |U  =�7   '  |�   >�7  |B  ?�7  |�  E�7   %'  |B   F�7  |C  G�7  |e  H�7  |8  I�7  |�  J�7  |

  X
8   0'  |�  Y
8  |�
  Z
8  }�   `38  ;'  |�  fD8   F'  |�  gD8  |�  hD8  |�  nm8   Q'  |�	  om8  |�  pm8  |H  v�8   \'  |`  w�8  |w  x�8  |   y�8  |~  �8   g'  |   ��8  |�  ��8  |  ��8  |�   ��8  |�  ��8  |�	  ��8  |�  �$9   r'  |  �$9  |  �$9  |�  �$9  |�  �Y9   }'  |�  �Y9  |�  �Y9  |�  �Y9  |m  ��9   �'  |	  ��9  |2	  ��9  |�  ��9  |9  ��9  |[  ��9   �'  |J  ��9  |�  ��9  |7  ��9  |�  �:   �'  |I	  �:  |$	  �:  |�   �-:   �'  |N  �-:  |p  �J:   �'  |�  �J:  |:  �J:  |�  �J:  |d   �J:  |�  ɋ:   �'  |  ʋ:  |�  ˋ:  |�	  Ѵ:   �'  |�  Ҵ:  |  ��:   �'  |�  ��:  |�  ��:  |�  ��:  |+  �;   �'  |�  �;  |�   �;  |  �/;   �'  |�
  �/;  |�  �/;  |  �X;   �'  |   �X;  |F  �X;  |�  �;   (  |�  �;  |�  ��;  |D  O�;   (  |�  P�;  |1  Q�;  |�  W�;    (  |^  X�;  |�  3�;   +(  |�  4�;  |�   8<   6(  |�  9<  |l	  =*<  A(  |N  >*<  |^  ?*<  |L  @*<  |a  D_<  L(  |B  E_<  |�	  F_<  |  G_<  |  H_<  |y  I_<  |�   �<   W(  |�  !�<  ~�� (  60  �DA0  �D�"%  �  �1  �<  (   �� O%  =  =  (  (   E=  �(    '   �_ � �� k  0M     � std  P  v  6�  x  K�  �  MP   x  Ob   m   R  P   	�  Qw  �   �   R   	�  R  �   �   R   
  T8  P  �   �   X   x  Z�   �   R   x  \�   �   R  ^   x  _�     R  �   x  c  #  R  i   �  p�  o  ;  F  R  ^   �  t�  o  ^  i  R  i   �  {y  �  R  u   n	 ~%  �  �  R  o   �  ��  |  �  �  X   �  �h  �  �  X    ;    :;   �  �d  � �  G�  c�� i�  �� .��   *     �� =�   %�  % �  J   �   ;   �  �  �  ;   ;   int �  �  �  '   �  !�� *   ")�  #  �)   ��  $ .  � %�)
   & � 0  P  #*  �)   �  %�)   & ?  P  '�  ['9  |"	 �   �a �� k� k  HM      std  ~  v  6�  x  K�  �  M~   x  Ob   m   �  ~   	�  Qw  �   �   �   	�  R  �   �   �   
  T8  ~  �   �   �   x  Z�   �   �   x  \�   �   �  �   x  _�     �  �   x  c  #  �  �   �  p�  �  ;  F  �  �   �  t�  �  ^  i  �  �   �  {y  �  �  �   n	 ~%  �  �  �  �   �  ��  �  �  �  �   �  �h  �  �  �    ;    :;   �  ��  � �  �� Dx  n  n   �� G%  +  �   �� �  @  K  �  �   (�  G� �  �  g  �    z �  ��  ;   �  �  �  ;   ;   int �  �  �  �  �  �  s  +  �  �   h  �   #  �   �  �  !K  �)   �  $  "h  $  �  �  #�  �� �)   �D  [  $�  � %�)&� �   #�  �� �)!   �v  �  $�  � '�  �)   �  (�  $� )�) *�)�   +�  �1  ~    ��   Jd �� g� k  �)�  � �  (  _� �>   �  int �  W   �  �  o  �	  �  qW  !E     "�   �  #  s  NL   �  VL   .  <z   `  DE   �  Wz   �  _�   �  eE   t   mE   a  uE     ~E   �  �E   3  �E   �  �E   H  �E   y  �E     �E   s  �E   T   �E   �  �E   F  �E   �  �E   �  �E     �E   V  �E   %   �  \	  2E   o  7E   �  <E   �  CE   �  E   �  �  %   `� �	    	$  
�  
3   
�    �� �O  3� �� � B� V�  <� �z  �� A� �� g� t�  �� �[  m�  �� O� �� �� /� �� ?� 5� k� 	p� 
�� O� +� �� J� �� �� �� M� � #� o� n� �� �� <� G� 8� �� �� �� ��  �� !+� "�� #�� $!� %{� &� 'f� (�� )�� *�� +�� ,~� -M� .� /'� 0�� 1�� 2�� 3�� 4�� 5� 6c� 7g� 8�� 9� :�� ;N� <�� =�� >J� ?�� � .� � o� � �� � � � [� � �� � ;� � �� � n� � �� � �� �  �}  s ��   len �E    ��  op ��    ]� 	%�  ,� 	(�   H�  	*�  len 	,E   Z}  	.E    �  �  ��  Z}  �E    H�  �%   �� �%  �� �z   u 0�   �  �\  �K  �%   B� �l   sat �l    ��  � �$   H�  �%   ��  � �O   H�  �%   �  ��     � 	M  H�  	P�   len 	RE   �� 	T�  @� 	VE   �� 	XC   
  �  
3  � �   len E    J  n� ,     a  �� E      �  < #%   � %%   (�  sub +%   num -E    �C  �� �[  u� �}  .� ��  �� �+  I� �\  a�  �  .� �  ��   �� 3  Q� J  >� &a  �� .�   �� 	3�  �  � � x� � � )� �� O� � 	 �� <	]I  s 	`�   ;� 	b�  �� 	dE   n 	f�  � 	h%  ]� 	jE   � 	lE   �� 	nI  �� 	pE    �� 	rE   $�� 	vE   (]� 	x%  ,~� 	|E   0�� 	~E   4p� 	�E   8 %  �� հ  ,� �%    w� ��  �� �E   '� ��  D� �E   �� ��  �� �E    �� ��  *5 ��   �� ��   �  �  �  �� �&	  *5 �&	   mod �  g� E    � �   �  �� 
n	  buf �   len 3   alc 3   $� E    �� �	  � �    � �   �� &�	  n (�   ]� )E   �� *E   �� +E   ~� ,E    /�	  W� � &� @0�
  buf 4�
   len 63    m� 9%   3� ;�  �� =�    � ?�  �� B&	  �� DE   m� GE   �� I>    � K   $ � ME   (� OE   ,2� Q�  0� SE   4.� UE   8�� W�  < %      �  � n	  �� Q%  -  di Q-  p S%   �  `� E   e  p %  s �  len E    W� E   �  p %  Z}  E   H�  %   �� ,E   �  p ,%  � -$  H�  .%   "� ?E     p ?%  � @O  H�  A%   �� �E     dc �%   l� 8,   _  di 8-   ��  :E    /� ;%   ret <,    �� %  �  di -  c E   p %   h� E   �  di -  c E    X� @%  �  di @-  i @,   p B%   �� �E     op �%   ,� ��   ]� �E   9  di �-  dc �%   �� `%  x  di `-  H�  `�  len `E   p b%   !K� s�  dpi s�   �	  �� yE   �  dpi y�   !� ��  dpi ��   k� �%   �  dpi ��   �� �%     Z}  �%  i �E   a �%   7� %  I  dpi �  dc �   *� �   }  dpi ��  � ��  i �E    !�� ��  dpi ��  s ��  l �3   i �3    !v� ��  dgs ��  � �3    �� �3    �� ��   ,	  �� P%  *  di P-  i P,   p R%   �� �%  _  di �-  ret �%   � �E    �� �%  �  di �-  �� �  p �%   !�� n�  di n-  �� n�   �	  !�� x�  di x-  �� x�    �%  2  di �-  �� �E    /� �%   "dc �%  "dcr �%     �� %  q  di -  num E   sub %  p %   � �%  �  di �-  op ��  p �%   !� �  dpi ��  �� �E   dc ��  �� �&	   � �E   " �� �E   p �&	    Y� UE   -  dc U�   �� WE    !�� cj  �� c�  �� cE   len c3   di d-   !u� ��  dgs ��  m� �3    !�� ��  dpi ��  �� �E   dc ��  �� �&	   �� �E    � �E   p �&	   �� �&	   !�� 48  dpi 4�  �� 4E   dc 5�  dpt 7�   !/� 'i  dpi '�  �� 'E   dc (�   6� �E   �  �� �E   dc ��  3� ��  �� ��   dpi ��	  " $� ��   �� ��    n	  �  #�   �  �  #�   (� �E   �  �� ��  �� �E   3� ��  �� ��   �Q  ��  �� �� ��   �� �/  di ��  dc �%   �� �E   " � ��   �� ��    �  �  #�   %  �  #�   �� ��    �� ��  �� �E   �� �  dgs �,	   �� �E    3   $z� _%  �)�   ��  %di _-  C� &�� _z  R&< `%  Q&� a%  � p c%  '  *hM �(  �� )hM *"  ��    $"� �%  �*F   �?  %di �-  �� +s ��  R+len �E   Qp �%  ,  �*   �  (  �� -�*   *"  ��   .3  �*    �(X  � (N  � (D  ��   /�� 
I  �*  ��  +di 
-  S&\ 
I  U&�� 
E   W v� 
I  0/� 
%   P)�M 1t 
z  R  $�� K
%  �+[   �4  %di K
-  )� %sub K
%  y� 2ret M
%  �� 3/� N
%   �� )�M 2t S
z  � 4.,  5Ps 5Q�R   $a� %  P,�  ��  %di -  G� 6P� E   �� 2c %   � 7�M �  3P� @E   q� 2p A�  �� 3w�  B�  �� 8�,   �  3/� G%   �  )�M 2s T�  2� 2len UE   P� 99  �,�M e[  (a  n� (U  �� (J  �� )�M :m  .  �-   d(  �� -�-   *"  ��     '9  s- N X(a  �� (U  �� (J  � ) N :m  '  s- N d(  � ) N *"  0�       )@N 2id s   C� )XN 3�� %s   ��    �  O  ;m� � .h   �\  6-� �\  �� 6�� �\  �� %dc ��  &� <M� +n.4w.�  5Pv 5Rw   E   !�� ��  dpi ��  c �%    =b  �.o   ��  (o  G� ({  � .�  �.;   �(�  ��   >   /t   �  ?/  �/  �*:  �� *F  �� *R  "�  $�� Y%  �/S   ��  %di Y-  _� ret [%  9  �/pN [c  (  _� )pN *"  ��   4�/�  5P�P#@/  �P  $�� I,   �/?   ��  %di I-  �� 2num K,   O� 4�/�  5Ps@/  s   $�� ]%   0U   �{  %di ]-  �� 3�� _,   �� 9�  G0�N jj  (�  � (�  .� )�N :�  .  G0   D(  .� -G0   *"  O�     4?0�  5Ps   $�� lE   �0#   ��  %di l-  b� 3�� n,   �� 4�0�  5P�P#@/  �P  �� g%    di g-  len gE    H�  i�  "s ��    $�� (%  �0�   �   %di (-  �� 2len *,   � ret +%  9�  �0�N 0�  (�  @� (�  t� )�N *�  �� 801@   �  *  �� 4h1�  5Ps 5R�4	5QE  A�0F�  4
1�  5Ps 5Rw 5Qv    4�0�  5Ps@/  s   >�  �1}   ��  (�  �� (�  � 8�1   ?  B�  ?�  S C�1�  [  5Pv @/  s  C�1�  w  5Pv @/  s  4�1�  5Ps@/  s   >   2q   �	  (1  T� ?=  �=  �9�  "2�N �  (  �� (�  �� )�N *  ��   .x  t2
   (�  �   $� &%  �2i   ��  %dpi &�  '� %dc '�  l� 2a )%  �� C�2	  d  5Pv  4�2�  5Pv 5Rs@=  �R  !�� ��  dgs ��  s ��  l �3    � �3    ;�� � 3�   ��  +s ��  � %l �3   �� 6�� ��   �� 2dgs ��  � '�  3�N �(�  N� ?�  � (�  � )�N *�  �� ,�  `3v   ��  (�  �� ?�  V-`3v   *�  �� *�  �� 8�3-   �  B�  ?�  V-�3-   :�  :�  A�3e�    A�3v�    AC3��     !�� ��  dpi ��  s ��   =�  �3�   ��  (�  � (�  @� ,}  �3|   ��  (�  l� (�  � (�  �� -�3|   *�  �� 'b  4O �({  �� (o  !� .�  :46   �(�  ?�     A�3��   !.� ��  dpi ��  l �,   buf ��   %   �  �   =�  �4�   ��   (�  R� (�  ~� D�  �G,�  �4�   ��   (�  �� (�  �� ,}  �4�   ��   (�  �� (�  �� (�  � -�4�   *�  4� 'b  �40O �({  S� (o  ~� .�  �4@   �(�  ��     A�4��   A�4��   !� �:!  dpi ��  H�  ��  len �E   p ��  end ��  "c �>   q ��  "dig �E      !�� x�!  dpi x�  � y�   �� {   src |�   �� |�!  "dst ��    �  E�� �@5�'  ��K  %dpi ��  �� 6�� �E   �� %dc ��  � 3�� ��  � 3� ��  p� 3-� �E   �� <F� lW7`O M$  2tp C  K� 9b  �5�O Tr"  ({  �� (o  �� .�  �U2   �(�  �   9b  �5�O V�"  ({  � (o  H� .�  �U2   �(�  q�   C�5�!  �"  5Ps 5Ru� C<6�!  �"  5Ps 5Ru� C�V�!  #  5Ps 5Ru� C�V�  $#  5Ps 5R	 C�V�  A#  5Ps 5R�	 C�Vb  [#  5Ps 5Rl C�Vb  u#  5Ps 5Ru C�V�  �#  5Ps 5R:6	 C�Wb  �#  5Ps 5R[ C�W�!  �#  5Ps 5Ru� C�Wb  �#  5Ps 5R] C�Wb  �#  5Ps 5R- C.\�  $  5Ps 5R�	 C�\b  3$  5Ps 5R- 4�\�  5Ps 5R�	  7�O �%  2sub 2�  �� ) P  �� 5   2a 6%  � 9I  H6HP 5�$  (Z  L� (Z  L� (f  u� )HP *r  ��   ,�  �6   M�$  (  � (�  %� -�6   *  %�   9:!  UR`P >s%  (S!  O� (G!  �� )`P *_!  �� *k!  �� *w!  �� 8�RO   [%  *�!  $   .x  �[   �B�     Cl6�  �%  5Ps  4�R�  5Ps    ,x  �6
   ��%  (�  M   7xP '  1len {E   W2i |E   n  2a }%  �  ,  �7   �&  (  �  -�7   *   �    ,�  �7d   ��&  B�  B�  .}  �7d   �B�  B�  B�  -�7d   *�   'b  �7�P �({  D (o  o .�  86   �(�  �      Cg7	  �&  5Ps  C�7�!  �&  5Ps 5Ru�5Qu� C�[w\  �&  5Ps 5Ru� 4�[�  5Ps 5RX6	  ,�  �8�   ��'  B�  B�  .}  �8�   �B�  B�  B�  -�8�   *�  � 'b  �8�P �({  � (o   .�  �8S   �(�  -      ,�  @9�   �6(  B�  B�  .}  @9�   �B�  B�  B�  -@9�   *�  @ 'b  @9�P �({  n (o  � .�  m9S   �(�  �      ,�  �9�   ��(  B�  B�  .}  �9�   �B�  B�  B�  -�9�   *�  � 'b  �9Q �({   (o  . .�  �9S   �(�  W      ,�  @:c   tT)  B�  B�  .}  @:c   �B�  B�  B�  -@:c   *�  j 'b  @:@Q �({  � (o  � .�  m:6   �(�  �      ,�  �:�   b6*  (�  
 (�  F -�:�   D�  ��,�  �:�   �+*  (�  Y (�  n '}  �:hQ �(�  � (�  � (�  � )hQ *�  � 'b  ;�Q �({  � (o   .�  =;S   �(�  5      A�:��    ,�  �;c   �*  B�  B�  .}  �;c   �B�  B�  B�  -�;c   *�  H 'b  �;�Q �({  v (o  � .�  �;6   �(�  �      9b  �;�Q p+  ({  � (o   .�  fU8   �(�  &   7�Q ]-  2op p%  9 3h� q%  � 3,� r�  ; 9b  �Q0R �+  ({  � (o  � .�  m[+   �(�  �   9b  �Q`R ��+  ({  � (o    .�  B[+   �(�     9b  SxR �,  ({  1 (o  S .�  �Z+   �(�  q   9b  ES�R �B,  ({  � (o  � .�  �Z+   �(�  �   Ct<8  d,  5Ps 5Ru�5Qw  C�<w\  �,  5Ps 5Ru�5Qu� C�Q8  �,  5Ps 5Ru�5Qu� C�Q�!  �,  5Ps 5Ru�5Qu� CES�Y   -  5Ps 5Ru�5Qu�#@   u� ClV�!  $-  5Ps 5Ru�5Qu� C�[w\  >-  5Ps 5Rw  4\8  5Ps 5Rw 5Qu�  ,�  �<c   f�-  B�  B�  .}  �<c   �B�  B�  B�  -�<c   *�  � 'b  �<�R �({  	 (o  0	 .�  �<6   �(�  Y	      7�R q/  2op R�  l	 2len SE   �	 ,�  0=�   U�.  (�  �	 (�  :
 .}  0=�   �(�  n
 (�  �	 (�  :
 -0=�   *�  �
 'b  0=S �({  �
 (o   .�  ]=S   �(�  J      ,}  �K   \3/  (�  ] B�  (�  � -�K   *�  � 'b  �K0S �({  � (o  � .�  L6   �(�  �     'b  �P�R X({   (o  % .�  6Z+   �(�  C    ,�  �=c   a 0  B�  B�  .}  �=c   �B�  B�  B�  -�=c   *�  V 'b  �=XS �({  � (o  � .�  �=6   �(�  �      7�S �0  2len 23   � 3�� 3>    ,�  `>d   8�0  B�  B�  .}  `>d   �B�  B�  B�  -`>d   *�   'b  `>�S �({  X (o  � .�  �>6   �(�  �      ,�  oS3   7�0  (�  �  4�M�!  5Ps 5Ru�  8�>;   �1  3�� E%  � 3�x F%  � C�>�!  81  5Ps 5Ru� C�>b  R1  5Ps 5R{ C�>�!  t1  5Ps 5Ru�5Qv  4�>b  5Ps 5R}  ,x  V?*   
�1  (�  �  ,�  �?c   f82  B�  B�  .}  �?c   �B�  B�  B�  -�?c   *�   'b  �?�S �({  9 (o  d .�  �?6   �(�  �      ,x  �?   �V2  (�  �  9�  @�S ��2  (�  � )�S *  �   7T 4  2op �%  	 3z  �%  6 3�� �%  X 3�� �%  � C9A�  �2  5Ps 5R56	 CNAw\  3  5Ps 5Ru�5Qu� CZAb  &3  5Ps 5R  CiA�!  H3  5Ps 5Rw 5Qu� CAw\  j3  5Ps 5Rw 5Qu� C�Zw\  �3  5Ps 5Rw 5Qu� C�Z8  �3  5Ps 5Rw 5Qu� C[w\  �3  5Ps 5Rw 5Qu� C[�  �3  5Ps 5R16	 4[w\  5Ps 5Rw 5Qu�  8�AW   f4  1dpm �  ��C�A�!  E4  5Ps 5Ru� 4�A�K  5Ps 5Ru�5Qu�  7 T K5  3�� �&	  � 0u� ��K  ��2i �s    3�� �&	  E ,x  �T   ��4  (�  y  C�B�!  �4  5Ps 5Ru� C�B�K  5  5Ps 5Ru� CCZU  25  5Ps 5Ru�5Qu�#@�  �Q 4Z�!  5Ps 5Ru�  7@T �7  2num �,   � ,�   Ef   ��5  B�  B�  .}   Ef   �B�  B�  B�  - Ef   *�  � 'b   E`T �({  � (o   .�  -E9   �(�  -      ,�   N_   ��6  B�  B�  .}   N_   �B�  B�  B�  - N_   *�  @ 'b   N�T �({  n (o  � .�  IN6   �(�  �      ,�  N�   �h7  (�  � (�  � -N�   D�  ��,�  �N�   �]7  (�   (�  4 .}  �Nu   �(�  R (�  � (�  � -�Nu   *�  � 'b  �N�T �({  � (o   .�  	O6   �(�  ,      A�N��    'b  ?O�T �({  ? (o  a .�  6X5   �(�      7�T H8  3H� ��  � 2a �%  � ,�  �S%   �8  (  � (�  � -�S%   *  �   CpE�  /8  5Ps 5Ru�#@=  u� 4�E�!  5Ps 5Ru�  7U W9  3� ^&	   2dcl _%  b 3�� `�  � C�E�!  �8  5Ps 5Ru� C	Fb  �8  5Ps 5R< CF�!  �8  5Ps 5Ru� C2Fb  �8  5Ps 5R> CpWb  9  5Ps 5R  C�Wb  !9  5Ps 5R  C�Y�!  =9  5Ps 5Ru� 4�Y�  5Ps 5Rl8	  ,}  RF�   �9  (�  � (�  
 (�   -RF�   *�  0 'b  pF0U �({  D (o  o .�  �FG   �(�  �     ,�  �Fc    f:  B�  B�  .}  �Fc   �B�  B�  B�  -�Fc   *�  � 'b  �FXU �({  � (o  � .�  G6   �(�  "      7�U �:  3b� �%  5 C�G�!  �:  5Ps 5Ru� CU�  �:  5Ps 5R�4	 CU�  �:  5Ps  4)U�  5Ps 5R�4	  ,}  �Gs   �f;  (�  k (�  � (�  � -�Gs   *�  � 'b  �G�U �({  � (o  � .�  �G6   �(�       7�U `<  3�� �&	  $ 3C� �%  k 0u� ��K  ��2i �s   � 1dpt ��  ��,x  �H   ��;  (�  �  7�U �;  3b� '%    CY�!  <  5Ps 5Ru� CCYb  +<  5Ps 5R  CPY�K  G<  5Ps 5Ru� 4�Y�!  5Ps 5Ru�  ,}  �Hx   ��<  (�  @ (�  f (�  y -�Hx   *�  � 'b  �H V �({  � (o  � .�  �H6   �(�  �     7(V 6=  1dpm o�  ��C�I�!  =  5Ps 5Ru� 4�M�K  5Ps 5Ru�5Qu�  7HV h=  3�� &	  � 4�S�!  5Ps 5Ru�  ,�  �Jc   ��=  B�  B�  .}  �Jc   �B�  B�  B�  -�Jc   *�  = 'b  �JhV �({  k (o  � .�  �J6   �(�  �      ,x  $K   �>  (�  �  9b  �L�V vV>  ({  � (o   .�  4U2   �(�  %   ,�   M_   ��>  (�  8 (�  P .}   M_   �(�  c (�  8 (�  P - M_   *�  w 'b   M�V �({  � (o  � .�  IM6   �(�  �      ,�  pOc   )�?  B�  B�  .}  pOc   �B�  B�  B�  -pOc   *�   'b  pO�V �({  ; (o  f .�  �O6   �(�  �      ,}  �O{   �@  (�  � (�  � (�  � -�O{   *�  � 'b   P�V �({  � (o  " .�  )P<   �(�  @     ,�  �Pg   �@  B�  B�  .}  �Pg   �B�  B�  B�  -�Pg   *�  S 'b  �P W �({  � (o  � .�  Q>   �(�  �      9�   THW ��A  (�   � (�   � (�    )HW *�   8 *	!  l 9b   TpW �A  ({  � (o  � .�  �T9   �(�  �   )�W *!  � * !  + 7�W HA  *+!  }  'b  H\�W �B{  (o  � .�  V\.   �(�  �      8V]   �A  1dpm ��  ��C:V�!  �A  5Ps 5Ru�	� 4ZVb  5Ps 5R   8aZ   +B  3ʗ ��  � ,x  iZ
   �B  (�  �  4�Zw\  5Ps 5Ru�  C�6�!  EB  5Ps 5Rv  C 7�  bB  5Ps 5R�6	 C7�!  |B  5Ps 5Rv  C7b  �B  5Ps 5R] C/7�!  �B  5Ps 5Rv  C;7�  �B  5Ps 5R�4	 CG7�!  �B  5Ps 5Rv  CS7b  C  5Ps 5R] C`8�  C  5Ps 5R�5	 Cp8�!  :C  5Ps 5Ru� C�8�  WC  5Ps 5R�6	 C�8�  kC  5Ps  C�8b  �C  5Ps 5R} C3<�!  �C  5Ps 5Rv  C?<�!  �C  5Ps 5Rv  C�<8  �C  5Ps 5Ru� C'>�!  �C  5Ps 5Ru� C+?�!  D  5Ps 5Ru� C7?b  'D  5Ps 5R  CQ?�  DD  5Ps 5R�5	 CK@w\  `D  5Ps 5Ru� C�@w\  |D  5Ps 5Ru� C�@b  �D  5Ps 5R) CaC�W  �D  5Ps 5Ru�	�5Qu�#@�  u� CyC�!  �D  5Ps 5Ru� C�C�  E  5Ps 5R35	 C�C�!  E  5Ps 5Ru� C�C�  ;E  5Ps 5R/5	 C�C�!  WE  5Ps 5Ru� C�C�  tE  5Ps 5R5	 C�C�!  �E  5Ps 5Ru� C�C�  �E  5Ps 5R5	 C�C�!  �E  5Ps 5Ru� CD�  �E  5Ps 5R�4	 CD�!  F  5Ps 5Ru� C/D�  F  5Ps 5R�4	 CAD�!  9F  5Ps 5Rv  CMD�  VF  5Ps 5R�4	 CYD�!  pF  5Ps 5Rv  CjD�  �F  5Ps 5R�4	 CzD�!  �F  5Ps 5Ru� C�D�  �F  5Ps 5R�4	 C�D�!  �F  5Ps 5Ru� C�Db  �F  5Ps 5R~ C�D�!  G  5Ps 5Ru� C�D�!  4G  5Ps 5Ru� CUG�!  NG  5Ps 5Rw  CkG�  kG  5Ps 5R�4	 C�I�  �G  5Ps 5R�5	 C�I�!  �G  5Ps 5Ru� C�I�  �G  5Ps 5Rp5	 C�I�!  �G  5Ps 5Ru� C
J�  �G  5Ps 5R`5	 CJ�!  H  5Ps 5Ru� C+J�  3H  5Ps 5RE5	 C;J�!  OH  5Ps 5Ru� CK�  lH  5Ps 5R�5	 CK�!  �H  5Ps 5Ru� CUKb  �H  5Ps 5R( C�K�!  �H  5Ps 5Ru� C�K�!  �H  5Ps 5Ru� C\L�Y  I  5Ps 5Ru�5Qw@   w  CnL�!   I  5Ps 5Ru� C�L�!  <I  5Ps 5Ru� C�L�!  XI  5Ps 5Ru� C�L�!  tI  5Ps 5Ru� C�L�  �I  5Ps 5R�6	 C�L�  �I  5Ps  C�Lb  �I  5Ps 5R} C	M�!  �I  5Ps 5Ru� C�M�!  �I  5Ps 5Ru� C�M�!  J  5Ps 5Ru� C�M�!  /J  5Ps 5Ru� C�Ob  IJ  5Ps 5R. C�P�W  qJ  5Ps 5Rv 5Qw@�  w  C�P�!  �J  5Ps 5Rv  C�W8  �J  5Ps 5Rw 5Qu� C�Wb  �J  5Ps 5R< C
X�!  �J  5Ps 5Rw  CX�  �J  5Ps 5R�6	 C%X�!  K  5Ps 5Rw  C1Xb  2K  5Ps 5R) C�Yb  LK  5Ps 5R[ C�Y�!  hK  5Ps 5Ru� C�Yb  �K  5Ps 5R] 41Z8  5Ps 5Ru�5Qu�  �  �K  �   E�� Z�\.  ��R  %dpi Z�  � 6�� ZE   k  %mod [�  �! 9b  �\�W l:L  ({  n# (o  �# .�  �b2   �(�  �#   ,�  @]p   ��L  B�  B�  .}  @]p   �B�  B�  B�  -@]p   *�  �# 'b  @]X �({  �# (o  $$ .�  q]?   �(�  X$      ,�  �]�   aXM  B�  B�  .}  �]�   �B�  B�  B�  -�]�   *�  k$ 'b  �]8X �({  �$ (o  �$ .�  ^O   �(�  �$      ,�  P^�   e�M  B�  B�  .}  P^�   �B�  B�  B�  -P^�   *�  �$ 'b  P^`X �({  "% (o  L% .�  �^O   �(�  j%      ,�  �^p   ivN  B�  B�  .}  �^p   �B�  B�  B�  -�^p   *�  }% 'b  �^�X �({  �% (o  �% .�  _?   �(�  �%      9b  @_�X v�N  ({  & (o  (& .�  c2   �(�  \&   9b  f_�X x�N  ({  z& (o  �& .�  �b2   �(�  �&   9b  �_�X {9O  ({  �& (o  �& .�  hc2   �(�  #'   ,�  �_p   }�O  B�  B�  .}  �_p   �B�  B�  B�  -�_p   *�  A' 'b  �_�X �({  {' (o  �' .�  �_C   �(�  �'      9b  I` Y rP  ({  �' (o  �' .�  �c2   �?�  S  ,�  �`�   ��P  B�  B�  .}  �`�   �B�  B�  B�  -�`�   *�  !( 'b  �`8Y �({  O( (o  y( .�  �`O   �(�  �(      ,�  0ap   �%Q  B�  B�  .}  0ap   �B�  B�  B�  -0ap   *�  �( 'b  0a`Y �({  �( (o  ) .�  aa?   �(�   )      9b  �a�Y �fQ  ({  3) (o  U) .�  �c2   �(�  ~)   ,�  �ap   �	R  (�  �) (�  �) .}  �ap   �(�  �) (�  �) (�  �) -�ap   *�  �) 'b  �a�Y �({  
* (o  4* .�  !b?   �(�  R*      9b  lb�Y �JR  ({  e* (o  �* .�  6c2   �(�  �*   F(]�!  C�a�!  mR  5Ps 5Rw  4lb�!  5Ps 5Rw   E�� � d�  �ZU  +dpi ��  V&�� �E   R&��  &	  S&�  E   U0H� �  W)�Y 0�� '&	  U1dc (%  S,�   eY   5S  B�  B�  .}   eY   �B�  B�  B�  - eY   :�  'b   e�Y �B{  Bo  .�  Je/   �B�       9b  ye Z 7�S  B{  Bo  .�  �eC   �B�    ,�  f]   =3T  B�  B�  .}  f]   �B�  B�  B�  -f]   :�  'b  f8Z �B{  Bo  .�  Ef3   �B�       9�  xf`Z >�T  B�  B�  )`Z D�  �G.�  �f�   �B�  B�  .}  �f�   �B�  B�  B�  -�f�   D�  U'b  �fxZ �B{  Bo  .�  �fB   �B�         .�  !gc   ?B�  B�  .}  !gc   �B�  B�  B�  -!gc   :�  'b  !g�Z �B{  Bo  .�  Lg8   �B�         =�  �g�  ��W  (�  �* (�  �* ?�  � ?�  ��  �*�  <+ 7�Z �V  *�  t+ *�  �+ ,�  �hp   FV  B�  B�  .}  �hp   �B�  B�  B�  -�hp   *�  �+ 'b  �h�Z �({  �+ (o  
, .�  �hB   �(�  (,      ,b  i^   �V  ({  ;, (o  P, .�  ,i4   �(�  c,   C�g�R  �V  5Ps 5Rv 5Q�  Ci�R  �V  5Ps 5Rv 5Q�  4j�R  5Ps 5Rv 5Q�   9b  �g[ &W  ({  v, (o  �, .�   j2   �?�  S  9b  �g0[ gW  ({  �, (o  �, '�  �iP[ �(�  -   9b  0hh[ !�W  ({  - (o  9- .�  `i@   �(�  e-   4*h�!  5Ps 5Rv   =�  `j&  ��Y  (�  x- (�  �- ?�  � ?�  ��  �*�  . *�  E. *�  �. *�  �. 9b  �j�[ �[X  ({  �. (o  �. .�  Tm2   �?�  S  9b  k�[ ��X  ({  / (o  L/ .�  k7   �(�  u/   9b  �k�[ ��X  ({  �/ (o  �/ '�  �l�[ �(�  �/   9b  �k\ �Y  ({  �/ (o  �/ .�  �l2   �(�  0   9b  bl(\ �_Y  ({  .0 (o  P0 .�  "m2   �(�  n0   Cxk�R  Y  5Ps 5Rw 5Qv  C�k�!  �Y  5Ps 5Rw  C�k�R  �Y  5Ps 5Rw 5Qv  4bl�R  5Ps 5Rw 5Qv   =�  �m5  ��[  (  �0 (  �0 ?   �   �D+  �h7H\ S[  B   (  !1 (  M1 )H\ :+  9b  #n`\ TzZ  ({  y1 (o  �1 .�  �n@   �(�  �1   9b  _n�\ Z�Z  ({  �1 (o  2 .�  �n@   �(�  K2   9b  o�\ S�Z  ({  ^2 (o  �2 .�  go/   �(�  �2   9b  @o�\ Y;[  ({  �2 (o  �2 .�  �o/   �?�  S  4Ln�!  5Ps 5Rw    C�m�!  m[  5Ps 5Rw  4�m�!  5Ps 5Rw   =8  �o�   �w\  (E  �2 (Q  63 (]  p3 8�oz   W\  (Q  �3 (]  �3 (E  �3 .}  �oq   +(�  4 (�  74 (�  J4 -�oq   *�  v4 'b   p�\ �({  �4 (o  �4 .�  )p7   �(�  �4      G�o�!  5P�P5R�R5Q�Q  E�� epp2  �y]  %dpi e�  �4 6�� eE   @5 %dc f�  v5 3}� hE   �5 9b  �p�\ o]  ({  6 (o  #6 .�  (qH   �(�  O6   9b  �p] rL]  ({  b6 (o  �6 .�  pq2   �?�  S  C�p�!  `]  5Pu  Gq�!  5P�P5R�X  �� t%  �]  di t-  �� tE   p v%   � �%  �]  di �-  �� �%   � ��   w�  ��  n �%   $�� �%  �q`  ��^  %di �-  �6 2ret �%  7 7(] �^  3�� �%  77 2t �z  v7 2s  �  �7 C�q�  y^  5Pv  CLr�  �^  5Pv  4[r  5Pv 5Ru 5Qw   'y]  �r@] �(�]  �7 (�]  �7 )@] *�]  �7 4�r�  5Pv 5R0    L� �%  _  di �-  ret �%   �� �%  `  di �-   /�  %   Ha_   �� 	%   H�  
%   Hs_   �U  E    H�_   H�  4%   H�_   �� G%   "op P%   ,� Q�   Z}  RE   H�_   h� w%   � xE    H�_   < �%   � �%   " z  �%   �� �%   �� �%     /�� p%  s�  �2g  +di p-  P X� r%  1al s%  �\1pal tI  S)X] a �%  '�^  `s�] �B_  )�] :_  '*  �s�] �B;  )�] :F  :R  '_  �s�] �B,_  )�] D7_  P7(^ �f  :�_  :�_  :�_  7x^ a  :�_  :�_   7�^ e  :�_  :`  D`  Q,_  �x)   �_a  B,_  -�x)   :7_  -�x)   :�_     9_  sy8_ ��b  B,_  )8_ D7_  P7�_ b  :�_  D�_  R:�_  7H` �a  :�_  :�_   7p` �a  D�_  VD`  WD`  P )�` :�_  D�_  V'�  ��` �B�  )�` D  P    7�` b  DH_  WDT_  V 8M}A   2b  :x_   7�` �b  Df_  Q.�  ~<   -B  B
  -~<   :  '  ~a TB  )a :"       )(a D�_  V   9_  *z@a ��c  B,_  )@a D7_  R7�a Ec  :�_  D�_  R:�_  7Hb �b  :�_  :�_   7pb c  D�_  VD`  WD`  P )�b :�_  D�_  V'�  @��b �B�  )�b D  P    7�b ]c  DH_  VDT_  W 8�}A   pc  :x_   7�b �c  Df_  Q.�  �~<   -B  B
  -�~<   :  '  �~c TB  )c :"       )(c D�_  V   '_  �z@c �B,_  )@c D7_  R7�c d  :�_  D�_  R:�_  7 d *d  :�_  :�_   7Hd Id  D�_  VD`  WD`  P )`d :�_  D�_  V'�  ���d �B�  )�d D  P    8�|L   �d  :x_   7�d �d  Df_  R.�  3   -B  B
  -3   :  .     TB  -   :"       7�d e  D�_  V )�d DH_  WDT_  V    )�d :�_  D�_  V9�  wpe �Re  B�  )pe D  P  '_  �{�e �B,_  )�e D7_  P7f �e  :�_  :�_  :�_  7Xf �e  :�_  :�_   7�f �e  D�_  WD`  VD`  P )�f D�_  VD�_  W'�  ��f �B�  )�f D  P    8�|F   	f  :x_   7�f if  Df_  P.�  �0   -B  B
  -�0   :  .  �   TB  -�   :"       7�f zf  D�_  V )�e DH_  WDT_  V     7g �f  Dx_  P 7 g g  Df_  R.�  �u.   -B  B
  -�u.   :  .  �u   TB  -�u   D"  Q     78g g  D�_  V )Pg DH_  WDT_  V         /� �%  ��  ��h  +di �-  U&� �%   R0�x �%  �\p �I  )pg arg �%  '*  ��g �B;  )�g :F  DR  P'_  ��g �B,_  )�g D7_  P7h [h  :�_  D�_  R:�_  7Hh h  :�_  :�_   7ph %h  D�_  VD`  WD`  P )�h :�_  D�_  V'�  "��h �B�  )�h D  P    7�h lh  Dx_  P 7�h �h  Df_  P.�  ��*   -B  B
  -��*   :  .  ��   TB  -��   D"  Q     7�h �h  D�_  V )i DH_  VDT_  W       $�� 	%   �#  �_�  %di 	-  8 3/� %   V8 2dim %  �8 9*  C� i �  (;  �8 ) i :F  *R  �8 '_  P�Pi �(,_  �8 )Pi *7_  �8 7xi �i  *�_  �9 C��2g  �i  5Ps 5RE Cј  �i  5Ps 5R05Qw  4מ�  5Ps   7�i V�  *�_  �9 *�_  �B *�_  2C 7�i @p  *�_  �C *�_  �C 9_  e��j ��o  (,_  �C )�j *7_  �D 7(k �m  *�_  �D *�_  yE *�_  F 7�k k  *�_  EF *�_  yF C�_  �j  5Ps  C�  �j  5Ps 5R55Qw  C׫_  �j  5Ps  C�  k  5Ps 5R7 4�2g  5Ps 5RE  7�k <l  *�_  �F *`  �F *`  G AC���  Cw�2g  _k  5Ps 5R_ C���  sk  5Ps  C��_  �k  5Ps  CΥ  �k  5Ps 5R:5Q�X C�  �k  5Ps 5R95Q�T C�  �k  5Ps 5R85Qw  C3�_  �k  5Ps  C>�_  l  5Ps  CI�_  %l  5Ps  4m�2g  5Ps 5RE  7�k {m  *�_  ^G *�_  �G 9�  )�l ��l  (�  H )l *  BH   CC�_  �l  5Ps  A\���  A|���  A����  C��J�  �l  5Ps  Cȧ  �l  5Ps 5R75Q�T C٧  m  5Ps 5R65Qw  C��2g  "m  5Ps 5RE C��  6m  5Ps  CU�_  Jm  5Ps  C�`  ^m  5Ps  4�  5Ps 5R45Q�X  C���  �m  5Ps  A����  C�  �m  5Ps 5R45Qw  4o��  5Ps   8�L   $n  *x_  zH C��J�  �m  5Ps  C�`  n  5Ps  4-�  5Ps 5R45Q�T  7 l �n  *f_  �H ,�  �0   -�n  (  �H (
  �H -�0   :  .  �   T(  �H -�   *"  �H     4q��  5Ps   78l o  *�_  I C��2g  �n  5Ps 5RE C��  �n  5Ps 5R05Qw  4a��  5Ps   7Pl �o  *H_  >I *T_  gI C���  6o  5Ps  C��J�  Jo  5Ps  CŪ  io  5Ps 5R15Qw  CӴ`  }o  5Ps  4�  5Ps 5R45Q�T  Cȡ_  �o  5Ps  Cۡ  �o  5Ps 5RI C���]  �o  5Ps  4���  5Ps    C�  p  5Ps 5R7 C1�  )p  5Ps 5R55Q�P 4��2g  5Ps 5RE  7hl J�  *�_  �I *`  �I *`  J 9_  J�Hm �v  (,_  :J )Hm *7_  JK 7�m �s  *�_  L *�_  lL *�_  �L 70n Gq  *�_  M *�_  HM C�_  �p  5Ps  C�  q  5Ps 5R55Qv  C�_  q  5Ps  C��  0q  5Ps 5R7 4V�2g  5Ps 5RE  7Xn jr  *�_  hM *`  �M *`  �M A���  C�2g  �q  5Ps 5R_ C��  �q  5Ps  CS�_  �q  5Ps  Ce�  �q  5Ps 5R:5Qw  Cx�  �q  5Ps 5R95Q�T C��  r  5Ps 5R85Qv  Cb�_  +r  5Ps  Cm�_  ?r  5Ps  Cv�_  Sr  5Ps  4�2g  5Ps 5RE  7�n �s  *�_  5N *�_  xN 9�  ѯ�n ��r  (�  �N )�n *  �N   C�_  �r  5Ps  A����  A���  A$���  C6�J�  �r  5Ps  CX�  s  5Ps 5R75Q�T Ci�  6s  5Ps 5R65Qv  C8�2g  Ps  5Ps 5RE C\��  ds  5Ps  Cl�_  xs  5Ps  CU�`  �s  5Ps  4g�  5Ps 5R45Qw   C���  �s  5Ps  A����  C��  �s  5Ps 5R45Qv  4���  5Ps   8$�F   Pt  *x_  #O C1�J�   t  5Ps  CN�`  4t  5Ps  4`�  5Ps 5R45Qw   7�n �t  *f_  AO ,�  ަ.   -�t  (  xO (
  �O -ަ.   :  .  ަ   T(  �O -ަ   *"  �O     4Ĩ�  5Ps   7�n 3u  *�_  �O C��2g  u  5Ps 5RE C
�  "u  5Ps 5R05Qv  4G��  5Ps   7�n �u  *H_  �O *T_  P Cγ�  bu  5Ps  C׳J�  vu  5Ps  C��  �u  5Ps 5R15Qw  C�`  �u  5Ps  4$�  5Ps 5R45Qv   C�_  �u  5Ps  C2�  �u  5Ps 5RI C���]  v  5Ps  4u��  5Ps    9_  �� o ��{  (,_  9P ) o *7_  �P 7�o �y  *�_  ,Q *�_  �Q *�_  KR 7p �v  *�_  �R *�_  �R C��_  �v  5Ps  C��  �v  5Ps 5R55Qv  C�_  �v  5Ps  C,�  �v  5Ps 5R7 4��2g  5Ps 5RE  7@p  x  *�_  �R *`  %S *`  gS A����  C��2g  Cw  5Ps 5R_ CƱ�  Ww  5Ps  C��_  kw  5Ps  C�  �w  5Ps 5R:5Q�X C#�  �w  5Ps 5R95Q�T C4�  �w  5Ps 5R85Qv  Cҹ_  �w  5Ps  Cݹ_  �w  5Ps  C�_  	x  5Ps  42�2g  5Ps 5RE  7hp _y  *�_  �S *�_  �S 9�  ���p �hx  (�  MT )�p *  �T   C�_  |x  5Ps  A'���  AG���  A_���  Cq�J�  �x  5Ps  C��  �x  5Ps 5R75Q�T C��  �x  5Ps 5R65Qv  C��2g  y  5Ps 5RE C���  y  5Ps  C��_  .y  5Ps  C��`  By  5Ps  4��  5Ps 5R45Q�X  CU��  sy  5Ps  CY�  �y  5Ps 5R45Qv  Aǲ��  4���  5Ps   8~�F   z  *x_  �T C��J�  �y  5Ps  C��`  �y  5Ps  4��  5Ps 5R45Qv   7�p �z  *f_  �T ,�  W�0   -|z  (  U (
  !U -W�0   :  .  W�   T(  !U -W�   *"  4U     4B��  5Ps   7�p �z  *�_  GU C°2g  �z  5Ps 5RE C԰  �z  5Ps 5R05Qv  4��  5Ps   7�p }{  *H_  }U *T_  �U C���  {  5Ps  C��J�  -{  5Ps  C��  L{  5Ps 5R15Qv  C�`  `{  5Ps  4��  5Ps 5R45Q�T  C��_  �{  5Ps  C��  �{  5Ps 5RI C���]  �{  5Ps  4���  5Ps    9_  ���p ���  (,_  �U )�p *7_  FV 7�q i  *�_  �V *�_  W *�_  �W 7�q �|  *�_  �W *�_  X C?�_  O|  5Ps  CS�  p|  5Ps 5R55Q�T C_�_  �|  5Ps  Cq�  �|  5Ps 5R7 4��2g  5Ps 5RE  7r �}  *�_  ?X *`  �X *`  �X Am���  C��2g  �|  5Ps 5R_ C���  }  5Ps  C�_  $}  5Ps  C��  E}  5Ps 5R:5Q�\ C�  f}  5Ps 5R95Q�X C�  �}  5Ps 5R85Q�T C&�_  �}  5Ps  C1�_  �}  5Ps  C<�_  �}  5Ps  4��2g  5Ps 5RE  70r   *�_  Y *�_  GY 9�  ��Pr �"~  (�  �Y )Pr *  �Y   C̭_  6~  5Ps  A���  A���  A���  C/�J�  e~  5Ps  CQ�  �~  5Ps 5R75Q�X Cd�  �~  5Ps 5R65Q�T C}�`  �~  5Ps  C��  �~  5Ps 5R45Q�\ C���  �~  5Ps  Cж_    5Ps  4+�2g  5Ps 5RE  C��  .  5Ps  A"���  CE�  X  5Ps 5R45Q�T 4H��  5Ps   8ΣL   �  *x_  Z CۣJ�  �  5Ps  C��`  �  5Ps  4�  5Ps 5R45Q�T  7hr J�  *f_  =Z ,�  �0   -9�  (  tZ (
  �Z -�0   :  .  �   T(  �Z -�   *"  �Z     4+��  5Ps   7�r ��  *�_  �Z C2�2g  v�  5Ps 5RE CF�  ��  5Ps 5R05Q�T 4x��  5Ps   7�r <�  *H_  �Z *T_  [ C���  ׀  5Ps  C��J�  �  5Ps  C��  �  5Ps 5R15Q�T C��`  �  5Ps  4�  5Ps 5R45Q�X  C_�_  P�  5Ps  Cr�  j�  5Ps 5RI C���]  ~�  5Ps  4���  5Ps    C>�2g  ��  5Ps 5R_ CG��  ��  5Ps  Cs�_  ҁ  5Ps  C��  �  5Ps 5R:5Qv  C��  �  5Ps 5R95Qw  C��  3�  5Ps 5R85Q�P 4��2g  5Ps 5RE  7�r �  *�_  8[ *�_  {[ 9�  B�`s ���  (�  �[ )`s *  �]   9_  T�xs �H�  (,_  z^ )xs *7_  S_ 7t $�  *�_  �_ *�_  �` *�_  �` 7�t u�  *�_  >a *�_  ra C�_  �  5Ps  C��  0�  5Ps 5R55Qv  C��_  D�  5Ps  C��  ^�  5Ps 5R7 4��2g  5Ps 5RE  7�t ��  *�_  �a *`  �a *`  b AN���  C~�2g  ��  5Ps 5R_ C���  Ѓ  5Ps  C��_  �  5Ps  Cϩ  �  5Ps 5R:5Qw  C�  %�  5Ps 5R95Q�X C�  E�  5Ps 5R85Qv  C�_  Y�  5Ps  C&�_  m�  5Ps  C/�_  ��  5Ps  4��2g  5Ps 5RE  7�t օ  *�_  Tb *�_  �b 9�  � u ���  (�  �b ) u *   c   C�_  �  5Ps  A���  A+���  A?���  CQ�J�  #�  5Ps  Cs�  D�  5Ps 5R75Q�X C��  d�  5Ps 5R65Qv  C�2g  ~�  5Ps 5RE CQ��  ��  5Ps  C�`  ��  5Ps  C�  Ņ  5Ps 5R45Qw  49�_  5Ps   C���  �  5Ps  A���  C��  �  5Ps 5R45Qv  4���  5Ps   8L�L   �  *x_  Xc CY�J�  N�  5Ps  Cx�`  b�  5Ps  4��  5Ps 5R45Q�X  7u �  *f_  wc ,�  �2   -��  (  �c (
  �c -�2   :  '  �0u T(  �c )0u *"  �c     4Ǥ�  5Ps   8R�=   b�  *�_  �c C_��  +�  5Ps  Cq�2g  E�  5Ps 5RE 4��  5Ps 5R05Qv   7Hu �  *H_  d *T_  /d C\��  ��  5Ps  Ce�J�  ��  5Ps  C��  ć  5Ps 5R15Qw  C˸`  ؇  5Ps  4ݸ  5Ps 5R45Qv   Cɢ_  �  5Ps  Cܢ  "�  5Ps 5RI Cۨ�]  6�  5Ps  4��  5Ps    CI�J�  \�  5Ps  Ck�  }�  5Ps 5R75Q�X C~�  ��  5Ps 5R65Q�P CC�2g  ��  5Ps 5RE C}��  ̈  5Ps  C��_  ��  5Ps  CX�`  �  5Ps  4j�  5Ps 5R45Qv   C-��  $�  5Ps  C�  E�  5Ps 5R45Q�P 4Ǟ�  5Ps   7`u ��  *x_  Xd CW�J�  |�  5Ps  C��`  ��  5Ps  4��  5Ps 5R45Qv   7xu 2�  *f_  �d ,�  ��.   -!�  (  �d (
  �d -��.   :  .  ��   T(  �d -��   *"  �d     4���  5Ps   7�u Ċ  *H_  �d *T_  e C��  a�  5Ps  C�J�  u�  5Ps  C-�  ��  5Ps 5R15Qv  C��`  ��  5Ps  4��  5Ps 5R45Qw   C��]  ؊  5Ps  C���  �  5Ps  C`�_   �  5Ps  4s�  5Ps 5RI     C�  .�  5Ps  C��  B�  5Ps  4��  5Ps 5R-5Qv   Y� �
%  |�  di �
-   � �
%  ��  di �
-   /� �
%   dim �
%  "s �
�    �� $%  �  di $-  cl &%  mem '%   $�� �%   �4  �	�  %di �-  7e 3/� �%   �e 2ret �%  �g 3�� �E   �g 9*  d��u �	.�  (;  �i )�u :F  *R  �j '_  n�(v �(,_  +k )(v *7_  �k 7�v �  *�_  �l *�_  �l *�_  Em 7�v Y�  *�_  �m *�_  �m C��_  �  5Ps  C�  �  5Ps 5R55Qv  C��_  (�  5Ps  C��  B�  5Ps 5R7 4��2g  5Ps 5RE  7w |�  *�_  �m *`  n *`  ^n A0���  Ca�2g  ��  5Ps 5R_ Cl��  ��  5Ps  C��_  ȍ  5Ps  C��  �  5Ps 5R:5Qu  C��  	�  5Ps 5R95Q�H C��  )�  5Ps 5R85Qv  C*�2g  C�  5Ps 5RE C��_  W�  5Ps  C��_  k�  5Ps  4��_  5Ps   70w ��  *�_  �n *�_  �n 9�  ��Pw �Ď  (�   o )Pw *  Io   C��_  ؎  5Ps  A����  A���  A(���  C:�J�  �  5Ps  C\�  (�  5Ps 5R75Q�H Cm�  H�  5Ps 5R65Qv  C��2g  b�  5Ps 5RE C��`  v�  5Ps  C�  ��  5Ps 5R45Qu  CY��  ��  5Ps  4i�_  5Ps   C»�  Ώ  5Ps  A����  C��  ��  5Ps 5R45Qv  4���  5Ps   8=�L   c�  *x_  �o CJ�J�  2�  5Ps  Ck�`  F�  5Ps  4�  5Ps 5R45Q�H  7hw �  *f_  �o ,�  H�2   -ؐ  (  �o (
  �o -H�2   :  .  H�   T(  �o -H�   *"  �o     4���  5Ps   7�w F�  *�_  p C��2g  �  5Ps 5RE C��  5�  5Ps 5R05Qv  4���  5Ps   7�w ؑ  *H_  Ep *T_  np Cy��  u�  5Ps  C��J�  ��  5Ps  C��  ��  5Ps 5R15Qv  C:�`  ��  5Ps  4L�  5Ps 5R45Qu   C��_  �  5Ps  C��  �  5Ps 5RI C���  �  5Ps  4���]  5Ps      7�w Ȓ  3\ �I  �p ,  ��   �n�  (-  �p ("  �p  8м    ��  2fn �%  �p  Cm�?  ��  5Ps 5R�\5Q0 C���  ��  5Ps  AżN�   ,   �$   �	�  (-  q ("  Iq  ,_�  P�   
	�  (p�  uq 4W�"�  5Ps   9|�  `��w 	��  (��  �q )�w *��  @r *��  �r 8��'   ��  :��  4���  5Ps 5Ru5Qv   9*  I�Px �
_�  (;  �r )Px :F  *R  ds '_  S��x �(,_  t )�x *7_  �t 7`y >�  *�_  \u *�_  �u *�_  Wv 7�y ��  *�_  �v *�_  �v C��_  *�  5Ps  C��  J�  5Ps 5R55Qw  CL�_  ^�  5Ps  C^�  x�  5Ps 5R7 4 �2g  5Ps 5RE  7�y ��  *�_  �v *`  1w *`  pw A����  C��2g  ֔  5Ps 5R_ C���  �  5Ps  C�_  ��  5Ps  C/�  �  5Ps 5R:5Qu  CB�  ?�  5Ps 5R95Q�H CS�  _�  5Ps 5R85Qw  C��_  s�  5Ps  C��_  ��  5Ps  C��_  ��  5Ps  4��2g  5Ps 5RE  7z �  *�_  �w *�_  �w 9�  ��0z ���  (�  >x )0z *  rx   C��_  �  5Ps  A����  A���  A*���  C<�J�  =�  5Ps  C^�  ^�  5Ps 5R75Q�H Co�  ~�  5Ps 5R65Qw  CP��  ��  5Ps  Ce�2g  ��  5Ps 5RE C��_  ��  5Ps  C�`  Ԗ  5Ps  4)�  5Ps 5R45Qu   C���  �  5Ps  A����  C��  -�  5Ps 5R45Qw  4	��  5Ps   7Hz ��  *x_  �x Cz�J�  d�  5Ps  C��`  x�  5Ps  4��  5Ps 5R45Qw   7`z �  *f_  �x ,�  �1   -	�  (  �x (
  y -�1   :  .  �   T(  y -�   *"  $y     4��  5Ps   7xz w�  *�_  7y Cw�2g  F�  5Ps 5RE C��  f�  5Ps 5R05Qw  4���  5Ps   7�z 	�  *H_  my *T_  �y C���  ��  5Ps  C��J�  ��  5Ps  C�  ٘  5Ps 5R15Qw  C�`  �  5Ps  4+�  5Ps 5R45Qu   C��_  �  5Ps  C��  7�  5Ps 5RI C���]  K�  5Ps  4��  5Ps      C��  s�  5Ps  4 �  5Ps 5R*5Qw    ,��  `�;   	�  (΋  �y -`�;   *ً  �y *�  �y Cm��  ݙ  5Ps  C~��  �  5Ps  4��  5Ps 5R+5Qv    7�z ��  3�� W	%   z ,_�  (�   i	V�  (p�  :z 4/�"�  5Ps   Cd�4  o�  5Ps 5R0 4{�`  5Ps   7�z H�  3Z}  A	%  Mz 3�� B	�	  kz ,�  �   D	К  (�  _{ (�  �{  ,�  7�    N	��  (�  �{ (�  �{  ,  ��%   H	�  (-  �{ ("  �{  C��  7�  5Ps 5R4 4+�`  5Ps   9_  ��z ���  ({  �{ (p  	| )�z :�  '  � { �(  	| ) { *"  |     9  R�{ :	ʛ  (-  /| ("  e|  ,_  ~�0   �	-�  ({  x| (p  �| -~�0   :�  .  ~�   �(  �| -~�   *"  �|     ,_  ��0   �	��  ({  �| (p  } -��0   :�  .  ��   �(  } -��   *"  }     ,_  ��0   �	�  ({  ,} (p  `} -��0   :�  .  ��   �(  `} -��   *"  s}     ,_  )�0   �	V�  ({  �} (p  �} -)�0   :�  .  )�   �(  �} -)�   *"  �}     ,_  n�0   �	��  ({  �} (p  ~ -n�0   :�  .  n�   �(  ~ -n�   *"  '~     ,_  ��0   �	�  ({  :~ (p  n~ -��0   :�  .  ��   �(  n~ -��   *"  �~     ,_  �0   �	�  ({  �~ (p  �~ -�0   :�  .  �   �(  �~ -�   *"  �~     ,  U�   �	��  (  �~ -U�   *"     C'�  ʞ  5Ps 5RA C��  ޞ  5Ps  C�  ��  5Ps 5R( Cͽ�  �  5Ps  C�  &�  5Ps 5R% C��N�  :�  5Ps  C��  N�  5Ps  C �  h�  5Ps 5R& C���  |�  5Ps  Cо  ��  5Ps 5R$ C��  ��  5Ps  C �  ğ  5Ps 5R" C��  ؟  5Ps  C0�  �  5Ps 5R# C��  �  5Ps  C���  �  5Ps  C̿  4�  5Ps 5R! C7��  H�  5Ps  Cy�`  \�  5Ps  Ci��h  p�  5Ps  C���  ��  5Ps  C��  ��  5Ps 5RI CP��  ��  5Ps 5R7	5Q4 C���  ܠ  5Ps@/  s  C���  �  5Ps  4���  5Ps@/  s   $�� �
%  `��   ���  %di �
-   1tl �
%  �\2ptl �
I  V )0{ 3�� �
%  � 3/� �
%   � C��  ��  5Ps 5R. 4���  5Ps    $�� �
%  @�d   �N�  %di �
-  � 6.� �
E   
� 32� �
%  (� 2tl �
%  Q� 3/� �
%   p� C\�	�  �  5Ps  Cr�  =�  5Ps 5R)5Qv  4���  5Ps   $�� i
%  ��[   ���  %di i
-  �� 2ret k
%  �� C����  ��  5Ps 5R1 4���  5Ps   �� %  �  di -  Z}  E   H�  	%  p %   $�� �%  ��  �ؤ  %di �-  /� 2c1 �%   e� 2c2 �%   �� 9��  i�H{ �ˣ  (٢  �� (͢  � (¢  E� )H{ :�  9  i�`{ ��  (  E� )`{ *"  Y�   'e  ~�x{ (�  l� (�  �� (v  Y�    7�{ n�  2low �E   �� 3�a  �E   ߂ )�{ 2i �E   �� 2p ��  G� 'q  $��{ (�  |� ?�  �\)�{ :�  .  ��   �?  �\-��   D"  P      8K�0   Ƥ  3�� �%  �� 3R� �E   �� Cb��  ��  5Ps  4x�  5Ps 5R3  4i�  5P�\  >� -%  �  di --  H�   � :$   " � VO    �� $%  T�  di $-  � $$  H�  %%  p '%   �� 2%  ��  di 2-  � 2O  H�  3%  p 5%   %� |%  ӥ  di |-  tl ~%  ret %  num �E    �� �%  �  di �-  ret �%  num �,    �� %  J�  di -  dc %   /� %   "tag 	%    $�� �%  ���  �B�  %di �-  ̃ 2ret �%  � 3/� �%   |� 9ӥ  +��{ -�  (�  � )�{ :�  *��  � ,  Q�   ���  (  3� -Q�   *"  F�   9  o��{ ��  (-  Y� ("  l�  4I��  5Ps    ,�  ��0   !��  ($�  � B�  -��0   */�  �� ) | *<�  �� C��  ��  5Ps  4��  5Ps 5RJ5Qu     ,��   ��   ]�  (��  ݅ - ��   *��  �� :��  *ƥ  � ,  L�   ��  (  -� -L�   *"  @�   9  u�| �7�  (-  S� ("  f�  C�	�  K�  5Ps  4D��  5Ps    9ؤ  ��0| ��  (�  y� 7P| �  *�  �� 'T�  ��p| n(|�  چ (p�  �� (e�  � )p| :��  9  ���| 7�  (  � )�| *"  +�   .�  ��6   8(�  >� (�  ]� (�  +�     - ��   *��  |� '�  ?��| Q(=�  �� (1�  އ (&�  �� )�| :I�  9  ?��| )��  (  �� )�| *"  �   .�  ]�3   *(�  #� (�  B� (�  �      C��  թ  5Ps  C���  �  5Ps  C��  ��  5Ps  C
�{  �  5Ps  CZ�  %�  5Ps  4l�  5Ps 5R55Qu    � o%  ��  di o-  ret q%   \ rI    � s%   N� �%  ߪ  di �-  ret �%  " /� �%    � �z  dc �%  " G� �%      `� 1%  "�  di 1-   H 3%  " H�  H%  num IE     $�� %  ���  ���  %di -  a� 3/�  %   �� 2dc !%  � 9ߪ  ���| )�  (�  �� )�| *��  ,� 7} ��  *�  v� *�  ̊ ,2  ��+   a�  (Z  � (N  $� (C  7� -��+   :f  .  ��   (  7� -��   *"  J�     C]�"�  0�  5Pv  C��  O�  5Pv 5R25Qs  C���  c�  5Pv  C��"�  w�  5Pv  C�{  ��  5Pv  4�{  5Pv   C��  ��  5Pv 5R0 C9�{  ɬ  5Pv  4R��  5Pv 5R7	5Q>   9B�  �(} &l�  (S�  ]� )(} D^�  �\*j�  �� *v�  � 9��  y�`} �5�  (��  � )`} *��  r� )h} *��  ӌ *��  � *Ī  b� ,  c�-   ���  (-  Í ("  ֍  7�} ǭ  *Ъ  � C���  ��  5Pv  A��J�   C7�J�  ۭ  5Pv  CQ�  ��  5Pv 5Qw  C��`  	�  5Pv  C�4  "�  5Pv 5R1 47��  5Pv     Co�?  T�  5Pv 5R�\5Q1 4���  5Pv 5Rw    ,  5�    a��  (-  	� ("  '�  7�} L�  3�� 0E   :� ,  	�'   OӮ  (-  Z� ("  m�  C�4  �  5Pv 5R0 C��`   �  5Pv  C��J�  �  5Pv  C���  6�  5Pv 5R(7	5Q3 4��  5Pv 5R1  C7�J�  `�  5Pv  C'�J�  t�  5Pv  C\�`  ��  5Pv  4��  5Pv 5R4  �� �%  �  di �-  H�   1� �%   ,� �,    �� �%   " H�  �%    �� %  R�  di -  p %   *5 %  len ,   i ,   c  %   str !�   .� �E   o�  dc �%   >�  ��$  ���  (�  �� (�  � *
  y� 7�} e�  (�  �� (�  �� )�} *
  N� )�} *  �� 9R�  ���} ��  Bc�  '  ��~ �(  ߐ   82�   �  *#  �  C��"�  3�  5Ps  C����  G�  5Ps  4��  5Ps 5R35Qv     '��  `� ~ �(��  � 9�  z�H~ ���  (�  G� )H~ *�  p� *�  ʑ *%�   � *1�  � *;�  y� *E�  Ȓ 9_  I�p~ G5�  ({  � (p  %� )p~ :�  .  I�   (  %� -I�   *"  C�     Ch��  I�  5Ps C���  i�  5Ps 5Rw 5Qv  C�  ��  5Ps 5R>5Q�\ 44�  5Ps 5R=5Q�\   8p�0   �  *�  V� Cw�"�  Ӳ  5Ps  C��  �  5Ps  4��  5Ps 5RF5Qv   8��P   }�  *��  t� *˯  �� *ׯ  �� C���  ?�  5Ps  C���  S�  5Ps C���  g�  5Ps  4��  5Ps 5R;  CG�"�  ��  5Ps  CZ�  ��  5Ps 5RC C���  ó  5Ps 5R0 C��  ܳ  5Ps 5RG C���  ��  5Ps 5R0 C�  �  5Ps 5RH C��  )�  5Ps 5Rv C+��  B�  5Ps 5R0 C>�  [�  5Ps 5R@ CM�"�  o�  5Ps  C`�  ��  5Ps 5RD Co��  ��  5Ps  C��  ��  5Ps 5R> C���  ϴ  5Ps 5Rh C���  �  5Ps 5R0 C
�  �  5Ps 5R? C��  �  5Ps 5R0 C,��  3�  5Ps 5R0 C=��  L�  5Ps 5R0 CP�  e�  5Ps 5RA C_�"�  y�  5Ps  Cr�  ��  5Ps 5RE C���  ��  5Ps  C��  ��  5Ps 5R9 C���  ӵ  5Ps  C��  �  5Ps 5R: C���   �  5Ps  C��  �  5Ps 5R= C���  -�  5Ps  C�  F�  5Ps 5RB C��  Z�  5Ps  C(�  s�  5Ps 5R< C���  ��  5Ps 5R0 4��  5Ps 5RG   >_  ��7  ��  (,_  Ó *7_  |� 7�~ �  *x_  �� C�J�  �  5Ps  C��`  �  5Ps  4��  5Ps 5R45Qv   7�~ X�  *�_  &� *�_  {� *�_  ߕ 7�~ ׷  *�_  .� *�_  b� C��_  r�  5Ps  C��  ��  5Ps 5R55Qu  Cw�2g  ��  5Ps 5RE C��_  ��  5Ps  4��  5Ps 5R7  7 ��  *�_  �� *�_  Ŗ 9�  ��0 ��  (�  � )0 *  C�   C��_  3�  5Ps  C�J�  G�  5Ps  C4�  h�  5Ps 5R75Q�X CE�  ��  5Ps 5R65Qu  C,�2g  ��  5Ps 5RE Ca��  ��  5Ps  C��_  ʸ  5Ps  C��`  ޸  5Ps  4��  5Ps 5R45Qv   7H �  *�_  {� *`  ŗ *`  � C;�2g  8�  5Ps 5R_ CD��  L�  5Ps  Cu�_  `�  5Ps  C��  ��  5Ps 5R:5Qw  C��  ��  5Ps 5R95Qv  C��  ��  5Ps 5R85Qu  C�_  Թ  5Ps  C�_  �  5Ps  C�_  ��  5Ps  4��2g  5Ps 5RE  Cf��  '�  5Ps  C[�  G�  5Ps 5R45Qu  4���  5Ps   7p ޺  *f_  P� ,�  ��:   -ͺ  (  |� (
  �� -��:   :  .  ��   T(  �� -��   *"  ��     4���  5Ps   7� ;�  *�_  �� Cl�2g  
�  5Ps 5RE C~�  *�  5Ps 5R05Qw  4���  5Ps   7� ͻ  *H_  � *T_  � C���  j�  5Ps  C�J�  ~�  5Ps  C&�  ��  5Ps 5R15Qv  Cu�`  ��  5Ps  4��  5Ps 5R45Qw   CA�_  �  5Ps  CT�  ��  5Ps 5RI F���]  F���   Q� �%  5�  di �-  s ��   !� Rr�  dpi R�  3� R�  �� S�   dc S�   =�  �D  ���  (�  H� (  f� (#  �� *Q  ؙ D]  ��|*h  � *s  W� I  9-  ��� ��  (^  j� (R  � (F  F� (:  f�  7� s�  J�  ��  �� J�  ��  :� 9�  I�8� ���  (*�  �� (�  	� Aw���  C���  q�  5Pw 5Ru�| 4O��  5Pw 5R0  ,i  ���   ���  (z  C� (�  W� (�  y� (�  �� -���   D�  ��}95�  ��X� �&�  (f�  �� (Z�  W� (N�  y� (B�  �� 4O��  5Pu`5RuT5Qv   7x� e�  J�  ��  � J�  ׿  � 4���!  5Ps 5RA5Qv   '�  ���� �(�  ,�    9y]  ��� �D�  (�]  [� (�]  {� )�� *�]  �� 9�]  ��Ѐ �-�  (�]  �� (�]  � )Ѐ *�]  � *�]  -� *�]  l� C���  �  5Pw  4��  5Pw 5RK5Qv    4M��  5Pw 5R1   C��  X�  5Pw  A����  4��  5P��|  K��  �� Kҿ  � K�  � A����   �  ��  L�  s�   �  %  ��  #�   n	  ҿ  L�  |�   �  �  �  L�  ��   �  MD� �  `�m  �%�  &�� �  � &z� �  �&�K    �&�� \  �3�� �  2� 2alc 3   [� 9�  ���� ) �  (�  �� (�  �� (�  � )�� D�  �P*�  � ,j  ��   ���  (�  M� (w  m�  C��r�  ��  5P� 5R 35Qt  A��e�    A����  A���  A�e�  Ai�e�   M�� jE   ��7   ���  &�� j�  � &3� k	  �&�� l�   �3�� nE   � 4��r�  5P� 5R�5Q�  ND  O��   �   N�  P��  N1  Q��  N�  W��   �   N^  X��  NU  =��   �   N�   >��  NB  ?��  N�  E�   �   NB   F�  NC  G�  Ne  H�  N8  I�  N�  J�  N

  Xd�   �   N�  Yd�  N�
  Zd�  O�   `��  �   N�  f��   �   N�  g��  N�  h��  N�  n��   �   N�	  o��  N�  p��  NH  v��   �   N`  w��  Nw  x��  N   y��  N~  %�     N   �%�  N�  �%�  N  �%�  N�   �%�  N�  �%�  N�	  �%�  N�  �~�     N  �~�  N  �~�  N�  �~�  N�  ���     N�  ���  N�  ���  N�  ���  Nm  ���   $  N	  ���  N2	  ���  N�  ���  N9  ���  N[  �)�   /  NJ  �)�  N�  �)�  N7  �)�  N�  �^�   :  NI	  �^�  N$	  �^�  N�   ���   E  NN  ���  Np  ���   P  N�  ���  N:  ���  N�  ¤�  Nd   ä�  N�  ���   [  N  ���  N�  ���  N�	  ��   f  N�  ��  N  �+�   q  N�  �+�  N�  �+�  N�  �+�  N+  �`�   |  N�  �`�  N�   �`�  N  ��   �  N�
  ��  N�  ��  N  ��   �  N   ��  NF  ��  N�  ���   �  N�  ���  N�  ���  N�  3�   �  N�  4�  N�   8!�   �  N�  9!�  Nl	  =>�  �  NN  >>�  N^  ?>�  NL  @>�  Na  Ds�  �  NB  Es�  N�	  Fs�  N  Gs�  N  Hs�  Ny  Is�  N�   ��   �  N�  !��  �  ��  �    0�� ���   2	��  �  �  �  = 0�� ��   .	��  O  /�  �   0<� �A�   -	�  P��  
9E   e�  
�  
�  
3    Q  ;v�  
�    P� R�   ��  
�   
3    R�d  �   ��  
�   
�  
�   PY2  
Q3   ��  
�   S�  6E   ��  
�  
�  T Uww  
BE   
�  
�    z	   �h (� �� �� �9  �; (  �  int �  �  L   �  �  o  �	  �  qW  !3     "�   �  #  s  NA   �  VA   .  <o   `  D3   �  Wo   �  _z   �  e3   t   m3   a  u3     ~3   �  �3   3  �3   �  �3   H  �3   y  �3     �3   s  �3   T   �3   �  �3   F  �3   �  �3   �  �3     �3   V  �3   �  \	  23   o  73   �  <3   �  C3   �  3   �� �3   � �h   �� ��   �� ��   �� �� �� p� �� �� �� �W  low ��   �a  ��   �v  	s �/  	ll ��   
�� �W  � ��  Y  n ��  d ��  rp �Y  nn �_  dd �_  rr �v  d0 ��  d1 ��  n0 ��  n1 ��  n2 ��  q0 ��  q1 ��  b ��  bm ��  ww �_  m1 ��  m0 ��    �  v  �� �  �9  �H  n �  � d �  ��  �� �   �  � �  � � �  �  � �  �  �� �  �� �  g� �  +� �  �� 
  ��   �    ,� *  צ 5  @� A  f� L  ��     D  OT   �   �  PT  1  QT  �  W}   �   ^  X}  U  =�   �   �   >�  B  ?�  �  E�   �   B   F�  C  G�  e  H�  8  I�  �  J�  

  X   �   �  Y  �
  Z  �   `9  �   �  fJ   �   �  gJ  �  hJ  �  ns   �   �	  os  �  ps  H  v�   �   `  w�  w  x�     y�  ~  �   �      ��  �  ��    ��  �   ��  �  ��  �	  ��  �  �*       �*    �*  �  �*  �  �_     �  �_  �  �_  �  �_  m  ��     	  ��  2	  ��  �  ��  9  ��  [  ��   "  J  ��  �  ��  7  ��  �  �
   -  I	  �
  $	  �
  �   �3   8  N  �3  p  �P   C  �  �P  :  �P  �  �P  d   �P  �  ɑ   N    ʑ  �  ˑ  �	  Ѻ   Y  �  Һ    ��   d  �  ��  �  ��  �  ��  +  �   o  �  �  �   �    �5   z  �
  �5  �  �5    �^   �     �^  F  �^  �  �   �  �  �  �  ��  �  3�   �  �  4�  �   8�   �  �  9�  l	  =�  �  N  >�  ^  ?�  L  @�  a  D	  �  B  E	  �	  F	    G	    H	  y  I	  �   l	   �  �  !l	   �	   j (� �� �� P�u  �< (  �  int �  �  L   �  �  o  �	  �  qW  !3     "�   �  #  s  NA   �  VA   .  <o   `  D3   �  Wo   �  _z   �  e3   t   m3   a  u3     ~3   �  �3   3  �3   �  �3   H  �3   y  �3     �3   s  �3   T   �3   �  �3   F  �3   �  �3   �  �3     �3   V  �3   �  \	  23   o  73   �  <3   �  C3   �  3   �� �3   � �h   �� ��   �� ��   �� �� �� p� �� �� �� �W  low ��   �a  ��   �v  	s �/  	ll ��   
�� �W  � ��  Y  n ��  d ��  rp �Y  nn �_  dd �_  rr �v  d0 ��  d1 ��  n0 ��  n1 ��  n2 ��  q0 ��  q1 ��  b ��  bm ��  ww �_  m1 ��  m0 ��    �  v  �� ��  P�u  �]  u ��  � v ��  �w ��  �� �  l�X� ��  �  �  �� �  L� X� �  �  �  �  .� �  �� �  C� �  �� �  �� 
  �   	�    5� *  z� 5  ��   A  �� L  ��     D  Oi   �   �  Pi  1  Qi  �  W�   �   ^  X�  U  =�   �   �   >�  B  ?�  �  E�   �   B   F�  C  G�  e  H�  8  I�  �  J�  

  X%   �   �  Y%  �
  Z%  �   `N  �   �  f_   �   �  g_  �  h_  �  n�   �   �	  o�  �  p�  H  v�   �   `  w�  w  x�     y�  ~  �   �      ��  �  ��    ��  �   ��  �  ��  �	  ��  �  �?       �?    �?  �  �?  �  �t     �  �t  �  �t  �  �t  m  ��     	  ��  2	  ��  �  ��  9  ��  [  ��   "  J  ��  �  ��  7  ��  �  �   -  I	  �  $	  �  �   �H   8  N  �H  p  �e   C  �  �e  :  �e  �  �e  d   �e  �  ɦ   N    ʦ  �  ˦  �	  ��   Y  �  ��    ��   d  �  ��  �  ��  �  ��  +  �!   o  �  �!  �   �!    �J   z  �
  �J  �  �J    �s   �     �s  F  �s  �  �   �  �  ��  �  ��  �  3�   �  �  4�  �   8�   �  �  9�  l	  =�  �  N  >�  ^  ?�  L  @�  a  D4	  �  B  E4	  �	  F4	    G4	    H4	  y  I4	  �   �	   �  �  !�	   �E   ~k � �� �� ���(  > (  _� �7   �  int �  �  W   �  �  o  �	  �  qW  !>     "�   �  #  s  NL   �  VL   .  <z   `  D>   �  Wz   �  _�   �  e>   t   m>   a  u>     ~>   �  �>   3  �>   �  �>   H  �>   y  �>     �>   s  �>   T   �>   �  �>   F  �>   �  �>   �  �>     �>   V  �>   �  \	  	2>   o  	7>   �  	<>   �  	C>   �  
>   �  �  E   	�� I  
��  
` 
�� 
j� 
�� 
� 
� 
� 
�� 
�  	
�� 

o� 
P 
J 
�� 
M  
� 
� 
� 
�� 
� 
�� 
h� 
� 
� 
�� 
�� 
Z� 
;� 
� 
�	 
�� 
�  
�� !
�� "
g #
� $
q� %
� &
'� '
�� (
�� )
�� *
1 +
�� ,
�  -
�� .
Y� /
�� 0
� 1
]� 2
*� 3
� 4
�� 5
)� 6
 7
� 8
 9
�� :
6	 ;
0 <
�� =
z� >
F� ?
�� � 
 � 
j  � 
� � 
Z� � 
b � 
� � 
� � 
 � 
#
 � 
�
 � 
  � 
� � 
 � 
�� � 

	 � 
z � 
�� � 
�� � 

 �  	� �D  
  
� 
�� 
O� 
0� 
�  	�� ��  
� 
�� 
o 
a 	
&� 

� 
�
 
�� 
�� 
�� 
� 
�� 
�� 
�� 
+	 
 
h	 
8 
3 
3� 
  
� 
� 
� 
�� 
�	 
��  
� !
� "
Z� #
D $
_ %
�� &
(� '
�	 (
�� )
�� *
h� +
S ,
r -
� .
@ /
M� 0
X� 1
c� 2
n� 3
y� 4
�� 5
�� 6
� 7
�� 8
�� 9
$ :
0 ;
< <
H =
T >
3� ?
� � 
N� � 
� � 
� � 
� � 
� � 
� � 
� � 
"� � 
� � 
� � 
� � 
	 � 
 � 
� � 
 � 
8
 � 
C
 � 
N
 � 
Y
 � 
d
 � 
o
 � 
z
 � 
� � 
�
 � 
�
 � 
�	 � 
D� � 
P� � 
\� � 
h� � 
t� � 
�	 � 
�� � 
�� � 
�	 � 
Q� � 
]� � 
i� � 
u� � 
� � 
�� � 
�� � 
�� � 
� � 
�� � 
T� � 
`� � 
c� � 
 � 
$ � 
�� � 
�� � 
I � 
U � 
a � 
m � 
y � 
< � 
I � 
V � 
c � 
� � 
.� � 
p �
} �
� �
� �
� �
� �
1  �
� �
� �
� �
� �
� �
� �
� �
� �
� �
\ �
I� �
G �
H� �
N �
-� �
�� �
� �
?� �
 �
�� �
C� �
�� �
& �
� �
�� �
�  �
� �
�
 �
< �
�� �
�� �
-� �
! �
7� �
�� �
 �
K �
�� �
�� �
�� �
� �
� �
.� �
U� �
�� �
o� �
�� �
�� � 	T ��	  
�� � 
%� �
>  �
  
�� 
� 
� 
� 
�	 
� 
H 
 
�� 	
s	 

M 
�� 
l 
2� 
 
�� 
N	 
� 
J� 
�� 
+� 
�
 
?� 
x� ?
�� 
�	 -
t .
 / + 0s     1>   (  5s   h  7s   �  =�   B6
  
�   
�  
M  
3  
�  
]  
K  
	  
�   �  L�	  �  WL
  R
  b
  6
  b
   h
  ^   Z�
  �  \�	   �  ]A
  V  b�	  `  c�	   �  n>   � ��
  �
  6
  �
  >   �
  �	  b
  �
  �    �
  �  ��g  reg �n   cfa ��   Hra ��   L  ��   P� �  Tn4 ��	  `�� ��	  d ��	  hA �~  l �� �r  x  6
  �  �
  �    � Ǘ  �  6
  �  >   �
  �	  b
  �
   �  %   2  7   �  �  l� �  �K  �P   � �E  P� ��   � UE  l� W�    � X�   ʗ Y�    �� j>   �� ks     nW   4� ��  �K  �P   � �E  �� �[  � ��  	 W   �  �   fde ��  )�  reg *�	  ,� +�	  exp ,�   �  W   .%  
�  
?� 
�� 
�� 
r� 
� 
6  (F  loc -�   how 6�   Aa  
��  
Y� 
�  � �&�  reg 7�   `  :�  �=� >�	  ��  ?�	  �� @�  �A� EF  � %  �  �   a  �"X  � Fa   pc I�   ��
 L�  � M�	  �i N�	  �� O�	  �� PW   ��� QW   �@� RW   �� SW   ��� T�   � { U�  
 n�   c  ~  �   E   �  �     ��  p ��   u2 �e   u4 �s   u8 ��   s2 �l   s4 �>   s8 ��    � pV  cfa �    �� �   =� %    %   \ V  �  e   X� e   Z�� ~  \ %   f  �   R�   ptr R�	  !&  R�	   N Rf  "� ��	  �  #�� ��
   $� ��  #�� ��
  %val �>    "�  ��	  �  #�� ��
   "j  ��  5  %p ��  %val �5  &�� �s   &  �W   &�T  ��   �  " 
 wc  W  %val w�	   '6 5�  (�� 5�
  (�U  5>   )p 5�    "  q�	  �  %val qc   *� *�   �  (�� *�
  (�U  *>    "K� ��   �  #�� ��
  #�U  �>    +� �	    (�� �
   +)  ��	  0  (�� ��
   +�  ��	  N  (�� ��
   +#  w�	  l  (�� w�
   "� ��   �  %p ��  ,up ��   �  �  "� �>   �  %p ��   "j �>   �  %p ��  ,up ��   "� �s   �  %p ��  ,up ��   "�
 �    %f ��     f  "� �<  <  %f �<   B  �  "� �>   a  %p ��   "�� �>   �  %p ��  ,up ��   "� �>   �  %p ��  ,up ��   "� �7   �  %p ��  ,up    "� �7   �  %p ��  ,up Ő   *B P>     (�� P�
  (�U  P>    -} *� ��	  B  (�� ��
   '�� �g  (�� ��
  )fs �g   X  .�  ��  ��A   ��  /p ��  ծ /val ��  � 0�� �s   � 0  �W   V� 0�T  ��  u�  �  *q  �    (�� �
  (�� W   )p �  )val    �	  "l  e�	  C  #�� eW   #�� e�
   "�  ��    #�� �W   #WC  ��	  %p ��  %val �    ��  ptr ��   u2 �e   u4 �s   u8 ��   s2 �l   s4 �>   s8 ��    ,u �  }  &�T  ��	  1�  ,a ��	   1
  ,tmp ��   2,tmp ��    �  3�� � ��	  �r  4 ��  �� 4r ��  � 4�� ��
  � 5fs �g  1� 6� ��  E� 7�  N��� ��  8�  �  9�� 6�  �W   � :reg ��  �� 6�� ��  #� 6,� ��  �� ;�� ��  �\7�  �ȁ �=  8  P� 8�  h� 9ȁ <  �� <  ڽ <)  �   =� �  >pc ��	  ?�  ��� �8	  /� 8�  g� 8�  �� 8�  /� 7  ��8� �  87  /� 8,  �� @0  1�	   t�  8A  [�  @N  ��   v�  8_  o�  A  ��   r8#  ��   ?C  :�`� 8r  �� 8i  ߿ 8^  �� 8S  �� 9`� <�  F� <�  ~� Bu�   �  C�  A�  u�   �D  8�  �� Eu�   <  �� <  � <)  2�    B��   �  F  �\G��m  HP�LHR��  E��   <�  P�      I�  ��   �.  D  8�  o� E��   <  �� <  �� <)  ��   I�  ��   �v  D  8�  �� E��   <  E� <  p� <)  ��   I�  ��0   ��  8  �� 8�  �� E��0   <  � <  :� <)  e�   I�  P�   �
  D  8�  �� EP�   <  �� <  �� <)  ��   I�  ��   R  D  8�  � E��   <  $� <  O� <)  b�   I�  ��   �  D  8�  u� E��   <  �� <  �� <)  ��   B�k   H  6T
 �  �� I�  �   �  D  8�  � E�   <  ^� <  �� <)  ��   J�  )�5   8  �� 8�  �� E)�5   <  � <  S� <)  f�    =�� b  6=� (�  ��  =�� |  6�� 8�  ��  I�  ��   @�  D  8�  �� E��   <  � <  D� <)  o�   7�  ���� B  8  �� 8�  �� 9�� <  �� <  � <)  <�   I�  P�   HT  D  8�  f� EP�   <  �� <  �� <)  ��   I�  ��   N�  D  8�  �� E��   <  � <  @� <)  S�   7�  ��Ђ V�  8  f� 8�  ~� 9Ђ <  �� <  �� <)  ��   I�  �   [,  D  8�  � E�   <  a� <  �� <)  ��   I�  @�+   bx  8  �� 8�  �� E@�+   <  � <  :� <)  M�   I�  ��   h�  D  8�  l� E��   <  �� <  �� <)  ��   I�  ��   t  D  8�  �� E��   <  � <  F� <)  |�   I�  `�   �P  D  8�  �� E`�   <  �� <  � <)  #�   I�  {�0   ��  8  B� 8�  Z� E{�0   <  �� <  �� <)  �   I�  ��   ��  D  8�  /� E��   <  ^� <  �� <)  ��   I�  @�   �,  D  8�  �� E@�   <  �� <  &� <)  9�   I�  p�+   �x  8  L� 8�  d� Ep�+   <  �� <  �� <)  ��   I�  ��   ��  D  8�  � E��   <  � <  D� <)  W�   I�  ��   �  8  v� 8�  �� E��   <  �� <  �� <)  �   K���E  L��m  +  HR�� L�m  A  HR�� L9�m  ^  HP�LHR�� G�m  HR��   *�� ��  �  )cie �  (�� ��
  )fs �g  >aug ��  >p ��  >ret ��  M�� ��  M�� ��  2M�
 ��	    "V  Hs      #�� HW    N� �6
   ��  �|&  4�� ��
  !� 5fs �g  r� :fde ��  �� :cie �  �� :aug ��  X� 6�  ��  �� :end ��  �� 7�  T�� ��   8�  i�  7r  �� � ��#  8�  �� D�  8�  �� 9 � <�  �� <�  � <�  �� <�  g� F�  �XI�  ��   �V!  D  8�  �� E��   <  �� <  �� <)  ��   I�  0�   ��!  D  8�  �� E0�   <  � <  2� <)  E�   =X� <#  C�  ?�  o��� �8	  X� 8�  �� 8�  q� 8�  �� 7C  o�Ѓ �"  8r  �� 8i  <� 8^  �� 8S  2� 9Ѓ <�  n� <�  2� =� Y"  F  �\G��m  HP�DHR�@  B��"   �"  C�  A�  ��"   �D  8�  �� E��"   <  �� <  �� <)  ��    E    <�  �    ?  �(� 87  �� 8,  q� @0  9�   t#  8A  :�  @       r #  8#  O�  AN  0    v8_  d�     Il  ��   �m#  8|  y� E��   <�  y�   I�  ��   ��#  D  8�  �� E��   <  �� <  �� <)  ��   K���E  G
�m  HR�X   I�  ��   ��#  8  ��  =P� �%  M  �	  ?�  p��� 8	  *� 8�  �� 8�  �� 8�  :� 7  p��� �$  87  :� 8,  �� @0  c�   tz$  8A  ��  @  �    r�$  8#  ��  AN  �    v8_  ��   ?C  ��Є 8r  �� 8i  
� 8^  �� 8S  � 9Є <�  I� <�  �� Bp�(   R%  C�  A�  p�(   �D  8�  � Ep�(   <  � <  B� <)  `�    B��   %  F  �\G��m  HPv HR�@  Bv    �%  <�  ~�  K���E      7"  �� � ��%  82  ��  7�  ��� ��%  8�  ��  =8� ;&  :i ��  k� J�   �   �D  8�  ~� E �   <  �� <  �� <)  ��    7"  1�P� Y&  82  ��  Kw��E  K��  GG�  HPw   OK� ��	  �&  #�� ��
  #�U  �>   &r �>   ,val �c   N� �	  � �  �;-  4�� �  �� 4  �  �� P�� �
  � P� �	  �;\y ;-  ��}6�� >   �� Q�� �P9h� :op D  �� 6�T  �	  �� :reg �  �� 6�� �  �� ;,� �  ��};�� �  ��}I�  p   a�'  8�  �� Ep   <�  ��   I|&  �=   �(  8�&  �� 8�&  �� E�=   <�&  �� <�&  �   =�� �)  Mj >�	  ?�  t�� ?8	  !� 8�  y� 8�  \� 8�  �� 7  t�� �(  87  �� 8,  \� @0  �   t�(  8A  �  @N  
   v�(  8_  *�  A  �   r8#  >�   ?C  � � 8r  R� 8i  �� 8^  �� 8S  �� 9 � <�  7� <�  � B�   :)  <�  W�  B   j)  F  ��}Gm  HP��}HR��}  EP   C�  A�  P   �D  8�  w� EP   <  �� <  �� <)  ��        7�  X� �*  D  8�  �� 9X� <  �� <  &� <)  E�   I|&  '>   �G*  8�&  X� 8�&  k� E'>   <�&  � <�&  ��   I|&  ~3   ��*  8�&  �� 8�&  �� E~3   <�&  �� <�&  ��   =p� �*  :t ��	  �  Ia  ?   ��*  8q  � E?   <z  �   =�� �*  6z  =�	  *� 6�� =�	  H�  =(� 4+  :t1 ��	  {� :t2 ��	  �� :t3 ��	  ��  I�  @    e|+  D  8�  �� E@    <  �� <  � <)  &�   I�  p   ��+  D  8�  9� Ep   <  Y� <  �� <)  ��   I|&  �3   �,  8�&  �� 8�&  �� E�3   <�&  �� <�&  ��   I�  `   !O,  D  8�  � E`   <  (� <  S� <)  f�   B�   �,  :ptr ��   y� Jl  �   �8|  y� E�   <�  y�    =@� �,  :ptr �   �� J�  %   8�  �� E%   <�  ��    K��E  L{m  -  HPw HR��} Lm  !-  HPw HR��} G�m  HPw HR��}   �	  K-  �  ? '� U�-  (�� U�
  )cfa U�   (�� V�-  Mr X>    �  '� @�-  (�� @�
  (�U  @>   )val A�	   3V� e��  �}2  4�� e�
  �� 5fs eg  A� ;� g�
  ��~:cfa h�   �� :i i%   �� ;�� {�  ��~I�  �   }X.  R�  8�  O�  IW  �   �.  8|  �� 8p  �� 8d  ��  B	B   /  :exp ��  � :len ��  ;� 7�  #	X� ��.  8  N� 8�  f� 9X� <  y� <  �� <)  ��   KZ	�&   7K-  �	p� ~o/  8p-  �� 8d-  �� 8X-  '� 9p� <|-  I� ?W  "�� a8|  {� Rp  Sd  ��~   I�-  �	   ��/  8�-  �� 8�-  �� 8�-  ��  7�  
�� ��/  8�  �� 8�  �  B@
[   �0  :exp ��  >� :len ��  h� >val ��	  I�  B
'   �K0  8  {� 8�  �� EB
'   <  �� <  �� <)  ��   IW  |
   �{0  8|    8p  "  8d  7   K|
�&   B�
p   H1  :exp ��  L  :len ��  v  :val ��	  �  I�  �
'   �1  8  �  8�  �  E�
'   <  �  <  �  <)     I�-  �
4   �>1  8�-  �  8�-  0 8�-  E  K�
�&   7W  �� �x1  8|  Z 8p  m 8d  �  I�      ��1  8�  � 8�  �  7W  @؇ ��1  8|  � 8p  � 8d  �  I|&  p@   �2  8�&   8�&  1 Ep@   <�&  G <�&  _   7�  ��� �s2  8�  � 8�  � T|&  �� �8�&  � 8�&  � 9 � <�&  � <�&  �    K�	�E   3* PD  ��3  4�� �
  > 4�� �   j 4�  �   � :ra �   � Ufs X  ��~;� �  ��~6,� 6
  � 7K-  �8� .i3  8p-  � 8d-  % 8X-  Q 98� <|-  } ?W  @X� a8|  � Rp  8d  �    V  �p   *L�   �3  HPv HRw  K��E  G�-  HPv HRw   3�� ��t   �i4  4�� ��
  � 5fs �g  F 7�  �x� �R4  8�  � 8�  � T|&  ��� �8�&  � 8�&  � 9�� <�&  � <�&   K��E     G��-  HPv HRw   Wc &6
   �   �C5  /exc &b
  q X�� '�
  � 0,� )6
   9�� Yfs -X  ��~0l� .>   E @$  �   35  85  } ?�  ��� �D�    L��3  5  HPv HRu  L�   85  HPv HRu  K��E    W� �6
  ��   �D6  /exc �b
  � X�� ��
   0� ��
  m 0{ ��   � 0,� �6
  � 0v� �6
  	 9�� Yfs �X  ��~0  �>   9	 @B  [	   �6  8[  q	 8O  �	 Gd�3  HPw HRu   Z(��~Lm   86  HPw HRu  Z���~  N� ^%   ��  �8  4I�  ^�
  �	 4\ _�
  
 :i a%   P
 ;� b�  �\I�  �   f�6  R�  8�  
  =� 7  :c k�   �
 :t l�   �
 98� :w q�	  ' >p r�	    7K-  6P� g{7  8p-  : 8d-  Z 8X-  z 9P� <|-  � 7W  Sp� ap7  8|  � 8p  � 8d  �  K;�E    7�  ��� ��7  8�  � 8�    E>'   6~� ��   d J�  >!   �8�  w 8�  � A|&  >!   �8�&  w 8�&  � E>!   <�&  � <�&  �      [|&  �X   �^8  S�&  � 8�&  � <�&   <�&  / K��E   [�  �   �z8  S  �  \$  �k   ��8  P�� �
  � 4�U  >   ^ ]val �	  �6r >   � :ptr �   � K'�E   ^�� Y�	  `   �9  P�� Y�
  �  ^  b�	  p   �d9  P�� b�
  � P�  bd9  �J�  x   dS�  �   >   \�  k�   ��9  P�� k�
  � ]val k�	  � ^�  q�   �   ��9  P�� q�
  �  [N  �   ��9  S_  �  ^� }�   �D   �6:  ]pc }�   � ;�   �d:fde ��   K��E   [0     �R:  SA  �  [      �n:  S#  �  ^6 %�:  0�   ��:  PY %�   � P�  %�:  �;�� '�
  ��}Ufs (X  ��~:reg )>   6 Gq   HPt HRw   �  3! C   �';  ]cfa C�   � P D�   � _�  R6
   c  �~<  /exc Rb
  I `$  T�
  ��|`>� T�
  ��}0,� U6
  � =�� �;  Yfs _X  ��~L��3  �;  HPu�|HRv  G�   HPu�|HRv   a$  ��� ��;  85  � J�  	   �D�    =Љ J<  0,� �%   � 0 ��    LJD6  @<  HP��|HR��| Ka�:   LM}2  d<  HPv HRu G4i4  HP� HR��|  b�� �6
  ��   �p=  /exc �b
  + X� İ
  c X{ Ğ   � `$  ��
  ��}`>� ��
  ��~0,� �6
  � =� >=  0,� �%   � 0 Ӟ    LD6  4=  HP��}HRw  K�:   L�}2  X=  HPv HRu G�C5  HPuHRw   cY  �@�   �b>  /exc �b
  # `$  ��
  ��}`>� ��
  ��~0,� �6
  [ = � >  0,� �%   y 0 �   � L�D6  >  HPu�}HRu�} K��:   Lx}2  *>  HPv HRu L�i4  G>  HPuHRu�} K��E  G�C5  HPu  b�  �6
   �   �N?  /exc �b
  � `$  ��
  ��}`>� ��
  ��~0,� �6
  � =� ?  6,� %    6 �   * L�D6  �>  HP��}HRw  K��:   LE}2   ?  HPv HRu L_C5  ;?  HPuHRw  Ki�E  K{';   d�� �   �t?  ]exc b
  �  e� 6
  ��   �2@  4 g  I 4p �   � ;�� �
  ��}6,� 6
  � =0� @  Ufs X  ��~LC�3  @  HPv HRu�} GP   HPv HRu�}  G}2  HPv HRu  fD  O>@   �   f�  P>@  f1  Q>@  f�  Wg@   �   f^  Xg@  fU  =�@   �   f�   >�@  fB  ?�@  f�  E�@   �   fB   F�@  fC  G�@  fe  H�@  f8  I�@  f�  J�@  f

  X�@   �   f�  Y�@  f�
  Z�@  g�   `#A  �   f�  f4A   �   f�  g4A  f�  h4A  f�  n]A   �   f�	  o]A  f�  p]A  fH  v�A   �   f`  w�A  fw  x�A  f   y�A  f~  �A     f   ��A  f�  ��A  f  ��A  f�   ��A  f�  ��A  f�	  ��A  f�  �B     f  �B  f  �B  f�  �B  f�  �IB     f�  �IB  f�  �IB  f�  �IB  fm  �~B   $  f	  �~B  f2	  �~B  f�  �~B  f9  �~B  f[  ��B   /  fJ  ��B  f�  ��B  f7  ��B  f�  ��B   :  fI	  ��B  f$	  ��B  f�   �C   E  fN  �C  fp  �:C   P  f�  �:C  f:  �:C  f�  �:C  fd   �:C  f�  �{C   [  f  �{C  f�  �{C  f�	  ѤC   f  f�  ҤC  f  ��C   q  f�  ��C  f�  ��C  f�  ��C  f+  ��C   |  f�  ��C  f�   ��C  f  �D   �  f�
  �D  f�  �D  f  �HD   �  f   �HD  fF  �HD  f�  �qD   �  f�  �qD  f�  �qD  f�  	3�D   �  f�  	4�D  f�   	8�D   �  f�  	9�D  fl	  	=�D  �  fN  	>�D  f^  	?�D  fL  	@�D  fa  	D	E  �  fB  	E	E  f�	  	F	E  f  	G	E  f  	H	E  fy  	I	E  f�  
 VE   �  f�  
!VE  W   wE  �   `� �gE  [hf� �iY2  Q,   �E  �   i� �<  �E  �   �E      D&   pq � � �� �  `L (  _� �7   �  int �  �  W   �  �  o  �	  �  qW  !>     "�   �  #  s  NL   �  VL   .  <z   `  D>   �  Wz   �  _�   �  e>   t   m>   a  u>     ~>   �  �>   3  �>   �  �>   H  �>   y  �>     �>   s  �>   T   �>   �  �>   F  �>   �  �>   �  �>     �>   V  �>   �  \	  2>   o  7>   �  <>   �  C>   �  	>   �  �  E   	�� 
I  
��  
` 
�� 
j� 
�� 
� 
� 
� 
�� 
�  	
�� 

o� 
P 
J 
�� 
M  
� 
� 
� 
�� 
� 
�� 
h� 
� 
� 
�� 
�� 
Z� 
;� 
� 
�	 
�� 
�  
�� !
�� "
g #
� $
q� %
� &
'� '
�� (
�� )
�� *
1 +
�� ,
�  -
�� .
Y� /
�� 0
� 1
]� 2
*� 3
� 4
�� 5
)� 6
 7
� 8
 9
�� :
6	 ;
0 <
�� =
z� >
F� ?
�� � 
 � 
j  � 
� � 
Z� � 
b � 
� � 
� � 
 � 
#
 � 
�
 � 
  � 
� � 
 � 
�� � 

	 � 
z � 
�� � 
�� � 

 �  	� 
�D  
  
� 
�� 
O� 
0� 
�  (  5s   h  7s   �  %   2  7   � !�  w #�   �� $,   t %�   �  �  �   �  �  l� ��  �K  �,   � �!  P� ��   -  �8 .�  t /  
 0$     �  r  4~  � 57    K 67     77    �� 87    �� ;7      3�  b <*  i =,    B� (�  P� *�    l� +�   � ,�   u 1�  s >~  *5 D�   �  � U!  l� W�    � X�   ʗ Y�    �� j>   �� ks    ls     nW   4� ��  �K  �,   � �!  �� �B  � ��  	 W   �  �   fde ��  ��  !>   | }�  �  >   �  �  �  �   �  �  � �  y �$   � �$   � �>   2  obj ��  f ��   G �>   N  �; �N   �  V 	>   r  �; 	N    � ��  7 ��  � ��   �  � d�    !ob d�  !pc d�   "vec f$  "lo g,   "hi g,   #"i k,   "f l  $P� m�   $� n7    �  j  �a  a  p �a  val �l  %�� �s   %  �W   %�T  �f   g  W   f  �
 ��  �  f ��   �  M  � ��  �  f ��   � =>   �  !f =�   &6 M	  S� M�  ob M�  l� N�   � N�    &� h'	  S� h�  ob h�   &m _	  S� �   ob �  l� ��   � ��    &? ��	  S� ��   ob ��   '' ݞ   �	  S� ��   (�  �a  �A   � 
  )p �a  � )val � 
   *�� �s   B *  �W   y *�T  �f  �  Z  +� J>   �   �m
  ,ob J�  � ,x K�  �,y K�  �-� MD  �#-� MD  �# .R ���   �  /ob ��  � 0+ ��  7 ,a �  � ,lo �>   �,hi �>   �1i �>   V 1j �>   � 2H�   1tmp ��  �  32�d3��d �  .�  ��   ��  /ob  �  � 0+  �  � 4� $  � 1a    1n 
,   ? 1m >   _ 2`� �  1tmp �  �  5m
  �  6P�h6R�l 7Bm
  6P�h6R�l  (V  Hs   `w   �	  8�� HW   � 9�	&   (k �D  �h   �I  8�� �W   D )ob ��  e 9	&   (�  �a  P/  ��  8�� �W   � 8WC  �D  � )p �a  � :val ��  �;  ��  ptr ��   u2 �e   u4 �s   u8 ��   s2 �l   s4 �>   s8 ��    <u ��  � �  *�T  �O  3 =�   B  <tmp �Z  �\7��	  6P� 6R�\  =     �  >tmp �f  ?       �@4  A+  } B     C?  � CJ  � CU  �    2x� �  Da �O  �  9U	&   D  �  +[ Y>   �{   ��  ,ob Y�  � ,x Y�  �,y Y�  �EWC  [D  & -� [D  �h-� [D  �l5�	  U  6Pv 6Ru  5�I  o  6Pv 6Rw  7�I  6Rw   + >      ��  /cie �  D 1aug 
a  � 1p 
a  � -R� D  �h$�� f  -�� Z  �lF  @	   2  @4  A+  } B@	   G?  CJ  � GU    F  `	   !r  @4  A+  � B`	   G?  CJ  � GU    F  p	   $�  A4  � A+  � Bp	   G?  CJ  � GU    9&  5T�	  �  6R�l 7�I  6R0  +� ^,   f  �*  /ob ^�  
 0� ^�  Z E� `�  � E�� a,   � E�� b>   L EWC  cD  � 2��   E g�   ErS  hD  B -P� hD  �lHr  [�� p�  A�  `  5o�  �  6Pw  5�	  �  6P�L6Ru  5�I  �  6P�L6R�T 7��  6P�L  I�     eA�  ~   . ��'  ��  /ob ��  � 07 ��  � 0� ��  � E� ��  � E�� �>   2 EWC  �D  [ 2؊ �  E ��  z 2 �   -P� �D  �lErS  �D  � 5T I  �  6P�X6R�P 7_ �  6P�X  =�   ,  1ptr �D  �  Fr  �   �S  A  � A�  �  Fr      �q  A�  �  5! �  �  6P�L 7- 	  6Ru   H�  � � ��  A�    7�	  6Pw 6Ru   J� �  � I  ��  ,ob �  P4� �  V,pc �   � $�  �  -�� !>   W$WC  "D  28� �  $ &�  -P� 'D  �h-� 'D  �l2h� �  $rS  DD  Kp Ea  P = !   �  $  <�   Ir  @!   1@�    I�   !   $@�    �  D  +, i>    "�   �B  ,ob i�  � ,x i�  �,y i�  �E k>   # E	 k>   6 -� lD  �h-� lD  �lH�  "�� n�  A�  I Fr  "   ?�  A�  I  9"�   H�  <"�� r�  A�  h Fr  <"   ?�  A�  h  9J"�   5*"	    6Pu 6R�  5<"I    6Pu  5X"	  1  6Pw 6R�  7i"I  6Pw    � ��  !ob ��  $7 ��  $�� �,   L� �M�  "p ��  #$� �,     M�  $� ��   #"p �    �  �  < �>   �  7 ��  �� �,   $r �,      ;6  !ob ;�  7 ;�  �� ;,   $+ =�    � ��  !ob ��  + ��  y �$  � �$  $/ ��  $�� �,   $a ��  "i �,   "j �,   "k �,   #$s ��       �  &  !ob  �  +  �  !v1 !$  !v2 !$  "i1 #,   "i2 #,   $� $�     ��  �  !ob ��  !pc ��   "vec �$  "lo �,   "hi �,   #"i �,   "f ��  $P� �D  $� �D  "p �a  $�� �>     � ~�  N  !ob ~�  !pc ~�   "vec �$  $�� �>   $WC  �D  "lo �,   "hi �,   #"i �,   "f ��  $P� �D  $� �D  "p �a    J� ��  �"n  �u  ,ob ��  U,pc ��   RH�  �"�� ��  @�  @�  N�� O�  VO�  UG�  N؋ G�  O�  PG�  G     HB  P#�� �Q  @O  N�� OZ  �XGf  Pr  �#=j#1   ,  O  VN(� O�  P  =�#   E  O�  4[ F�  J%S   u  @�  @�  BJ%S   O�  V  2@� �  O�  V Q�  �%X� @  @  @  NX� O)  WH6  -&�� J  @f  @Z  @N  @C  N�� G~  G�  G�  G�  G�  Or  0[N�� G�     I�  p(�   M@�  @�  @�  @�  Bp(�   G  G  G        =�#O   �  Kp ��  VB�#   Kf ��  P  H&  @$Ќ �  @B  @7  NЌ GM  GY  Gd  N� Gp  Oz  WO�  �TO�  �XO�  PG�  Q�  �$� �@�  Ir  �$   ?@�       Q�  �& � �@�  @�  N � G�  G�  G�  O�  QG
  N8� G  O   VO*  �TO6  �XOB  P    R�   *V   ��  A�  � A�  � A�  � A�  � B*6   A�   A�  $ A�  D A�  c   R	  `*W   ��  A	  � A	  � S�  s*   j2  T�   T�   A�  � A�  �  B�*7   A	    A	     ?�  �*7   j@�  @�  @�  @�  B�*7   T�   T�   A�    A�         U� n�*c   �j  VS� n�   � Dob p�  @  S	  �*9   w`  A	  @  A	  S  B�*9   A	  @  A	  S  ?�  �*9   j@�  @�  @�  @�  B�*9   A�  f  A�  f  A�  @  A�  S      9�*%&   R'	  0+K   ��  A3	  z  A>	  �  AH	  �  AS	  �   R_	  �+K   ��  Ak	  ! Av	  /! W'	  �+X� �TS	   TH	   A>	  N! A3	  !   U\ ��+V   �  VS� ��   � <ob ��  PS_	  �+;   �u  Xv	  PAk	  m! ?'	  �+;   �TS	   TH	   X>	  PA3	  m!   9�+%&   Y� ��   0,�   ��  8S� ��  �! Dp ��  �! Dob ��  +" Zout �9�,	&  9-:&   �  R�	   -   �  X�	  � [%-  6� �   U� �0-2   �c  VS� �   � S�	  I-	   �Y  A�	  �" 9R-   9Z-:&   \� ��  p-   ��   ,pc ��   � 4� ��   �1ob ��  �" 1f ��  �" L& =�-Z   [   E�� >   ## -ʗ D  �\F�  �-   0   A�  e# Fr  �-   ?&   A�  e#  9�-�   5�-	  J   6Pw 6Rv  7
.I  6Pw   2p� �   1p ��  x# 7U.N  6Pu 6Rw   7�-N  6Pv 6Rw   �  ]D  O�    �   ]�  P�   ]1  Q�   ]�  W�    �   ]^  X�   ]U  =�    �   ]�   >�   ]B  ?�   ]�  E!!   �   ]B   F!!  ]C  G!!  ]e  H!!  ]8  I!!  ]�  J!!  ]

  Xn!   �   ]�  Yn!  ]�
  Zn!  ^�   `�!  �   ]�  f�!   �   ]�  g�!  ]�  h�!  ]�  n�!   �   ]�	  o�!  ]�  p�!  ]H  v�!   �   ]`  w�!  ]w  x�!  ]   y�!  ]~  /"     ]   �/"  ]�  �/"  ]  �/"  ]�   �/"  ]�  �/"  ]�	  �/"  ]�  ��"     ]  ��"  ]  ��"  ]�  ��"  ]�  ��"     ]�  ��"  ]�  ��"  ]�  ��"  ]m  ��"   $  ]	  ��"  ]2	  ��"  ]�  ��"  ]9  ��"  ][  �3#   /  ]J  �3#  ]�  �3#  ]7  �3#  ]�  �h#   :  ]I	  �h#  ]$	  �h#  ]�   ��#   E  ]N  ��#  ]p  ��#   P  ]�  ��#  ]:  ��#  ]�  ®#  ]d   î#  ]�  ��#   [  ]  ��#  ]�  ��#  ]�	  �$   f  ]�  �$  ]  �5$   q  ]�  �5$  ]�  �5$  ]�  �5$  ]+  �j$   |  ]�  �j$  ]�   �j$  ]  �$   �  ]�
  �$  ]�  �$  ]  �$   �  ]   �$  ]F  �$  ]�  ��$   �  ]�  ��$  ]�  ��$  ]�  3%   �  ]�  4%  ]�   8+%   �  ]�  9+%  ]l	  =H%  �  ]N  >H%  ]^  ?H%  ]L  @H%  ]a  D}%  �  ]B  E}%  ]�	  F}%  ]  G}%  ]  H}%  ]y  I}%  ]�  	 �%   �  ]�  	!�%  _ ,�  @[_ -�  <[]" 0�   `f� �aY2  Q,   %&  �   a�� E�   :&  ,    b  ;�     %U  $ >   :;I  $ >      I  :;n   :;I8  	 :;I8  
9:;   :;  .?:;I<   I     & I  &   I  .?:;I<  .?:;I<  .?:;<  . ?:;I<  .?:;<  .?:;n@�B   :;I  ���B1  �� �B  4 :;I  4 :;I  .?:;<   %U  $ >   :;I  $ >      I  :;n   :;I8  	 :;I8  
9:;   :;   <  & I  <  .?:;2<d   I4  . ?:;n<  .?:;I<   I     &   I  .?:;I<  .?:;I<  .?:;<  . ?:;I<  .?:;<  9:;  :;  .:;I<  .:;I<   4 :;I<  !. ?:;I<  ".?:;n<  #. ?:;<  $.?:;n<  % :;  &:;n  '(   (  ) <  * :;I  +: :;  ,.G   - :;I  . :;I  /.:;   0 :;I  1  24 :;I  3.:;I   44 :;I  5.:;I   6 I  7.G d  8 I4  9.:;I@�B  : :;I  ;  <4 :;I  =.:;I@�B  > :;I  ?4 :;I  @ :;I  AU  B4 :;I  C  D4 :;I  E��1  F�� �B  G4 :;I  H1XY  I 1  J 1  K4 1  L�� 1  M:;  N :;I  O :;I  PU  Q1RUXY  R :;I  S1XY  T 1  U��1  V.G@�B  W :;I  X
 :;  Y
 :;  Z4 :;I  [4 :;I  \4 :;I  ]1RUXY  ^1XY  _4 1  `1RUXY  a1XY  b:;  c:;  d.4<d  e.:; d  f.:; d  g4 :;I  h4 :;I  i4 :;I  j4 G  k. ?:;<  l.?I4<  m. ?4<  n.?4<  o.?n4<   %U  9:;   :;I  .?:;nI@�B   :;I  �� 1     $ >  	.?:;nI<  
 I  .?n4<  .?4<   %U  9:;  9:;  :;   :;I8  .?:;<cd   I4   I  	.?:;n<d  
.?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   :;   :;I   <  . ?:;nI<  . ?:;n<      I   I  ;   B I  $ >  $ >  :;n   :;I8   :;I   :;n  !(   "  #:;  $ :;I8  %.:;I<  &.:;I<  '.?:;<  (. ?:;<  )4 :;I<  *.?:;n<  +.?:;<  ,. ?:;I<  -.?:;I<  . :;  /   0: :;  1.G   2 :;I  3.:;   4 :;I  5  64 :;I  7 :;I  8.1@�B  9 1  :U  ;4 1  <�� 1  =U  > 1  ?�� �B1  @.G@�B  A :;I  B :;I  C  D4 :;I  E1XY  F4 G  G.?:;I<  H.?:;I<   %U  $ >   :;I  $ >      I  :;n   :;I8  	 :;I8  
9:;   :;   <  . ?:;n<  .?:;I<   I     & I  &   I  .?:;I<  .?:;I<  .?:;<  . ?:;I<  .?:;<  :;n  (     :;  9:;  .:;I<  .:;I<   4 :;I<  !.?:;n<  ".?:;I<  # :;  $: :;  %.G   & :;I  ' :;I  (.?:;@�B  ) :;I  *1XY  + 1  ,  -4 :;I  .�� 1  /4 :;I  04 :;I  14 G   %U  $ >   :;I  $ >   I     &   & I  	 :;n  
9:;   :;   :;  9 :;  :;  .?4<d   I4  / I  /   /   .?:;n<   I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   :;I8  .?:;2<d  .?:;nI2<d  .?:;n2<d   I82    :;I2  !.?:;2<d  ":;  # I8  $ :;I8  %.?:;<d  &.?4<d  ' :;I?2<  ( :;I?<  ). ?:;nI<  *.?:;nI<d  +.?:;n<d  ,.?:;n<d  -.?:;nI<d  ..?:;nI<d  /.?:;n<  0. ?:;nI<  1.?:;2<d  2.?:;2<cd  3.?:;nI2<d  4.?:;nI2<d  5.?:;n2<d  6.?:;nI<  7/ I  8 <  9 :;I?2<  : :;I?2<  ;:;2  < :;I?<  =.?:;n<d  ><  ?.?:;2<cd  @:;2  A.?:;<d  B.?:;2<d  C.?:;nI2<d  D.?:;nI2<  E. ?:;nI2<  F.?:;<cd  G. ?:;n<  H:;  I(   J :;I2  K :;I?2<  L :;I?2<  M :;I?2<  N:;  O I8L2  P I842  Q.?:;L2<d  R.?:;nI2<d  S.?:;L2<d  T.?:;n2<d  U.?:;nILM2<d  V<  W.?:;I<  X.?:;<  Y.?:;I<  Z :;I?2<  [. ?:;n<  \9:;  ]/ I  ^.:;I<  _.:;I<  `: :;  a I  b. ?:;I<  cI  d!   eI  f   g I  h.G   i :;I  j  k4 :;I  l.G d  m I4  n :;I  o4 :;I  p :;I  q4 :;I  r :;I  s. G   t.G:; d  u.G:; d  v.1n@d�B  w 1  x 1  y1XY  z�� �B  {1XY  |1RUXY  }��   ~�� �B1  ���B1  ��� �B  ��� 1  �.G@d�B  � I4  � :;I  ����B�B  �.G@d�B  �.1n@d�B  �  �4 1  �1XY  �U  �4 1  �1RUXY  �1RUXY  �U  �4 :;I  �4 I  �4 :;I  � 1  � 1  � :;I  �4 :;I  �4 :;I  �1RUXY  �1XY  � 1  �4 1  � :;I  �  �.G@�B  �.G@�B  �.1n@�B  � :;I  � :;I  � :;I  � I4  �4 :;I  �4 :;I  �.?n4<  �. ?4<  �.?I4<  �.?nI4<   %U  9:;  9 :;   :;  :;   :;I  .?:;n<   I  	& I  
.?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   :;I8  .?:;2<d   I4  .?:;nI2<d  .?:;n2<d  / I   I82   :;I2  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I?<  . ?:;nI<  .?:;nI<d   .?:;n<d  !.?:;n<d  ".?:;nI<d  #.?:;nI<d  $.?:;n<  %. ?:;nI<  &.?:;2<d  '.?:;2<cd  (.?:;nI2<d  ).?:;nI2<d  *.?:;n2<d  +.?:;nI<  ,/ I  - <  .:;  /(   0<  1 :;I2  2 :;I?2<  3 :;I?2<  4 :;I?2<  5.?:;L2<d  6.?:;nILM2<d  7.?:;n<d  8.?:;I<  9. ?:;n<  :9:;  ;/ I  <:;  =.?:;nILM2<d  >.?L42<d  ?$ >  @$ >  A: :;  B :;I  C I  D   EI  F&   G  H :;n  I I  J. ?:;I<  KI  L!   M.?:;<  N.?:;I<  O. ?:;I<  P.?:;<  Q.G d  R I4  S.G:; d  T.G   U :;I  V :;I  W. G   X :;I  Y  Z4 :;I  [ :;I  \.1n@d�B  ] 1  ^ 1  _1XY  `�� �B  a1XY  b��   c�� �B1  d.G@d�B  e I4  f�� 1  g  h4 :;I  i :;I  jU  k4 :;I  l4 :;I  m I4  n4 1  o4 1  p 1  q4 :;I  rU  s1RUXY  t4 1  u.G@d�B  v :;I  w1RUXY  x 1  y.G@�B  z :;I  {1XY  |1XY  }.G@�B  ~1RUXY   1  �1RUXY  �4 :;I  �.?:;I<   %U  $ >   :;I  $ >   I     &   & I  	 :;n  
9:;   :;  9 :;  :;  .?:;n<   I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I8    :;I?<  !. ?:;nI<  ".?:;nI<d  #.?:;n<d  $.?:;n<d  %.?:;nI<d  &.?:;nI<d  '.?:;n<  (. ?:;nI<  ).?:;2<d  *.?:;2<cd  +.?:;nI2<d  ,.?:;nI2<d  -.?:;n2<d  ..?:;nI2<d  /.?:;nI<  0/ I  1/ I  2 <  3 :;I?2<  4 :;I?2<  5:;2  6 :;I?<  7.?:;<d  8.?:;n<d  9:;2  :.?:;<d  ;.?:;2<d  <.?:;nI2<d  =.?:;nI2<  >. ?:;nI2<  ?.?:;<cd  @. ?:;n<  A:;  B(   C<  D :;I2  E :;I?2<  F :;I?2<  G :;I?2<  H :;I?<  I :;I?<  J.?:;nI2<d  K.?:;nI2<d  L.?:;n2<d  M.?:;n2<d  N.?:;I<  O/ I  P.?:;nI<  Q9:;  R: :;  S I  T. ?:;I<  UI  V!   W.G d  X I4  Y :;I  Z :;I  [  \4 :;I  ].G   ^ :;I  _4 :;I  ` :;I  a. G   b4 :;I  c.G@d�B  d I4  e :;I  f :;I  g :;I  hU  i4 :;I  j4 :;I  k4 :;I  l1XY  m 1  n1RUXY  o  p4 1  q1XY  r  s�� 1  t1RUXY  uU  v4 1  w1RUXY  x 1  y1RUXY  z1XY  {4 I  |��   }.G@�B  ~1XY   :;I  � :;I  �4 :;I  �4 :;I  �4 :;I  �4 :;I  � 1  � 1  �4 1  �4 :;I  �4 :;I  �4 :;I  �.?nI4<  �.?I4<  �. ?4<  �.?n4<   %U  $ >   :;I  :;   :;I8   I  9:;   :;  	 :;  
 I8  9 :;  / I  /   /   .?:;n<   I  & I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   :;I8  .?:;<d  .?4<d    :;I?2<  ! :;I?<  ". ?:;nI<  #.?:;nI<d  $.?:;n<d  %.?:;n<d  &.?:;nI<d  '.?:;nI<d  (.?:;n<  ). ?:;nI<  *.?:;2<d  +.?:;2<cd  ,.?:;nI2<d  -.?:;nI2<d  ..?:;n2<d  /.?:;nI2<d  0.?:;nI<  1/ I  2 <  3 :;I?2<  4 :;I?2<  5:;2  6 :;I?<  7.?:;n<d  8<  9.?:;2<cd  :.?:;n2<  ;. ?:;nI2<  <.?:;nI2<  =:;2  >.?:;<d  ?.?:;2<d  @.?:;nI2<d  A.?:;nI2<  B.?:;<cd  C. ?:;n<  D :;I?<  E :;I?<  F:;  G(   H :;I2  I :;I?2<  J :;I?2<  K :;I?2<  L:;  M:;2  N.?:;n2<  O:;2  P(   Q.?42<d  R:;2  S:;2  T :;I  U:;  V :;I?2<  W.?:;L2<d  X.?:;nILM2<d  Y0 I  Z:;  [.?:;L<d  \ :;I82  ].?:;I2<d  ^:;  _ :;I82  `.?:;n2<d  a:;  b.?:;<d  c.?:;L<d  d.?:;nLM2<d  e/ I  f.?:;I<  g.?:;nI2<d  h   i. ?:;n<  j.?:;n<  k$ >  l. ?:;I<  m I  n   o&   p :;n  q9:;  r.:;I<  s.?:;I<  t.?:;I<  u: :;  v I  wI  x!   y:;  z! I/  {.G   | :;I  }  ~4 :;I  .G d  � I4  �4 :;I  � :;I  � :;I  � :;I  �4 :;I  �.G:; d  �.G:; d  �. G   �4 :;I  �   �.4   �.1n@d�B  � 1  ����B  ��� �B  �.G@d�B  � I4  �.G:;@d�B  � I  � :;I  �U  �4 :;I  �1XY  ���   ��� 1  ��� �B  ��� �B1  �1XY  � 1  ����B1  �.1n@d�B  �.1@d�B  �1RUXY  � 1  �1RUXY  �4 1  � :;I  �U  �4 :;I  �4 :;I  �1RUXY  �1XY  �1RUXY  ���1  �1XY  �.1@d�B  �4 :;I  � 1  �  �  �.G@�B  � :;I  � :;I  �.1n@d  �4 1  �4 1  �.G@d�B  � :;I  � :;I  �4 :;I  ��� �B  �4 1  �4 :;I  �4 :;I  � 1  �4 :;I  �.G@�B  � 1  �4 :;I  �4 :;I  �.4@�B  �4 :;I  �4 :;I  �4 Gn  �.?I4<  �.?n4<  �.?nI4<  �. ?4<  � <  �. ?I4<  �.?nI4<   %U  9:;  9 :;   :;   :;I  :;   I82  .?:;2<d  	 I4  
 I  .?:;2<d  & I  4 :;nI?<  9:;   :;   :;I2  .?:;nI2<d  .?:;n2<d  / I  $ >  $ >  : :;   I  &    I  .G d   I4  .1n@d�B   1   :;I  .1n@d�B   %U  $ >   :;I  :;   :;I8   I  9:;   :;  	9 :;  
.?:;n<   I  & I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I?<  . ?:;nI<  .?:;nI<d  .?:;n<d   .?:;n<d  !.?:;nI<d  ".?:;nI<d  #.?:;n<  $. ?:;nI<  %.?:;2<d  &.?:;2<cd  '.?:;nI2<d  (.?:;nI2<d  ).?:;n2<d  *.?:;nI2<d  +.?:;nI<  ,/ I  -/ I  . <  / :;I?2<  0 :;I?2<  1:;2  2 :;I?<  3.?:;<d  4.?:;n<d  5<  6.?:;n2<  7:;2  8.?:;<d  9.?:;2<d  :.?:;nI2<d  ;.?:;nI2<  <. ?:;nI2<  =.?:;<cd  >. ?:;n<  ? :;I?<  @ :;I?<  A:;  B :;I82  C :;I82  D :;I?2<  E :;I?2<  F :;I2  G.?:;2<cd  H.?:;nI2<d  I.?:;L2<d  J.?:;nILM2<d  K.?:;n<d  L.?:;I<  M$ >  N. ?:;I<  O   P&   Q :;n  R9:;  S.?:;n2<d  T/ I  U:;  V: :;  W I  XI  Y!   Z:;  [:;n  \ :;I8  ]   ^I  _.?:;I<  `.?:;I<  a.?:;<  b.?:;<  c! I/  d.G d  e I4  f.4   g :;I  h.G@d�B  i I4  j :;I  k :;I  l.1n@d�B  m 1  n�� 1  o�� �B  p��   q�� �B1  r :;I  s.G@d�B  t I4  uU  v4 :;I  wU  x4 :;I  y1XY  z 1  {4 :;I  |1XY  }4 :;I  ~4 :;I  4 Gn  �.?n4<  �.?I4<  �.?nI4<   %U  $ >   :;I  $ >   :;I   I     :;  	 :;I8  
I   I  &   & I     :;n  9:;   :;  9 :;  .?:;n<  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;  (   <  :;2   :;I?<  .?:;2<d   I4  .?:;2<d    :;I2  !.?:;nI2<d  " :;I2  #.?:;nI2<  $ :;I?2<  % :;I?2<  & :;I?2<  '.?:;2<cd  (/ I  )/ I  *.?:;nI2<d  +.?:;L2<d  ,.?:;n2<d  -: :;  ..?:;nI2<d  /.?:;L2<d  0.?:;n2<d  1.?:;I<  2.?:;nI2<d  34 :;nI?<  44 :;nI?<  59:;  6.:;I<  7.:;<  8.?L42<d  9<  : I  ;. ?:;I<  <.?:;<  =.?:;I<  >. ?:;I<  ?.?:;<  @.G   A :;I  B  C4 :;I  D.G d  E I4  F :;I  G4 :;I  H.G:; d  I :;I  J. G   K.?:;I   L :;I  M.?:;   N.1@�B  O 1  P1RUXY  Q 1  R 1  S1XY  T��   U1RUXY  V1XY  W�� 1  X  Y4 1  Z1XY  [.1n@d�B  \ 1  ]U  ^4 1  _���B1  `�� 1�B  a 1  b�� �B1  c.G@�B  d :;I  eU  f4 :;I  g4 :;I  h��1  i4 :;I  j4 :;I  k4 :;I?<  l.?n4<  m.?I4<  n. ?4<   %U  9:;   :;  :;   I8  9 :;   :;   :;I  	:;  
 I82  .?:;2<d   I4   I  .?:;2<d  & I   :;  9  4 :;I<  : :;  9:;  4 :;I<  :;  0 I  :;   <  .?:;n<  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   (   !<  " :;I2  # :;I2  $ :;I?2<  % :;I?2<  & :;I?2<  '.?:;nI2<d  (.?:;n2<d  ).?:;L2<d  */ I  +/ I  , :;I8  -.?:;nI2<d  ..?:;nI2<d  /.?:;nI2<d  0.?:;n2<d  1.?:;I<  24 :;nI?<  39:;  4.?:;n2<d  5/ I  6:;  7 :;I  8 :;I8  95 I  :.?:;<d  ;.?:;n<d  <.?:;nI<d  = :;I  >.?:;nI<d  ?.?:;n<  @.?:;2<d  A :;  B :;I8  C <  D:;  E :;I?2<  F :;I?<  G.?:;nI2<  H.?:;n2<  I.?:;nI2<d  J4 :;I<  K: :;  L:;  M$ >  N$ >  O   P :;I  Q I  R:;n  S :;I8  T   U&   VI  W.?:;I<  X.?:;I<  Y.?:;<  Z. ?:;I<  [.?:;<  \ I  ]  ^ :;n  _I  `! I/  a. ?:;I<  b.G d  c I4  d :;I  e.G   f :;I  g. G   h :;I  i.1n@d�B  j 1  k1RUXY  l 1  m�� �B  n1XY  o��   p�� 1  q�� �B1  r.G:;@�B  s :;I  tU  u4 :;I  vU  w4 :;I  x  y4 :;I  z  {4 :;I  | :;I  }4 1  ~4 1  1XY  �1XY  �.G@d�B  � I4  �4 :;I  �4 :;I  �4 G  �4 G  �4 G:;n  �.?n4<  �.?:;n<   %U  $ >   :;I  $ >   I  & I   :;n  9:;  	 :;  
9 :;  :;  .?:;n<   I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  <  .?:;nI2<d   I4   :;I2  .?:;n2<d  / I  / I  .?:;nI<   :;I8  .?:;I<  . ?:;I<  9:;  : :;   I   .G d  ! I4  " :;I  #.G   $  %4 :;I  & :;I  '. G   (.G@�B  ) :;I  *U  +4 :;I  ,4 :;I  -1RUXY  . 1  /  04 1  11XY  2 1  34 1  41XY  51XY  64 1  71RUXY  8  91RUXY  : 1  ;1RUXY  <4 :;I  =4 :;I   %U  $ >   :;I  $ >   I     &   & I  	 :;n  
9:;   :;   :;  :;   I8  9 :;  .?:;n<   I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   :;I8  .?:;2<d   I4  .?:;nI2<d  .?:;n2<d  / I   I82   :;I2  .?:;2<d   :;  ! :;I8  ".?:;<d  #.?4<d  $ :;I?2<  % :;I?<  &. ?:;nI<  '.?:;nI<d  (.?:;n<d  ).?:;n<d  *.?:;nI<d  +.?:;nI<d  ,.?:;n<  -. ?:;nI<  ..?:;2<d  /.?:;2<cd  0.?:;nI2<d  1.?:;nI2<d  2.?:;n2<d  3.?:;nI<  4/ I  5 <  6:;  7(   8<  9 :;I2  : :;I?2<  ; :;I?2<  < :;I?2<  =.?:;L2<d  >:;  ? :;I82  @.?:;nI2<d  A.?:;n2<d  B.?:;nILM2<d  C.?L42<d  D:;  E.?:;2<cd  F.?:;L2<d  G.?:;n2<d  H.?:;n2<d  I.?:;I<  J/ I  K.?:;I<  L9:;  M:;  N :;I82  O.:;I<  P: :;  Q I  R. ?:;I<  SI  T!   U.G   V :;I  W  X4 :;I  Y.G d  Z I4  [ :;I  \4 :;I  ] :;I  ^ :;I  _. G   `.G:; d  a   b.G@d�B  c I4  d  e4 :;I  f1XY  g 1  h4 1  i1RUXY  jU  k :;I  l  m1XY  n 1  o1RUXY  p.1@d�B  q 1  r�� 1  s.G:; d  t.1n@d�B  u 1  v1RUXY  w1XY  x1RUXY  y��   zU  {4 1  |1XY  }��1  ~�� �B   :;I  � :;I  � I4  � :;I  � :;I  � 1  �4 :;I  �4 :;I  � :;I  �4 1  � :;I  �4 :;I  �4 :;I  �.?n4<   %U  $ >   :;I  $ >   I     &   & I  	 :;n  
9:;   :;  9 :;  :;  .?:;n<   I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I8    :;I?<  !. ?:;nI<  ".?:;nI<d  #.?:;n<d  $.?:;n<d  %.?:;nI<d  &.?:;nI<d  '.?:;n<  (. ?:;nI<  ).?:;2<d  *.?:;2<cd  +.?:;nI2<d  ,.?:;nI2<d  -.?:;n2<d  ..?:;nI2<d  /.?:;nI<  0/ I  1/ I  2 <  3 :;I?2<  4 :;I?2<  5:;2  6 :;I?<  7.?:;<d  8.?:;n<d  9:;2  :.?:;<d  ;.?:;2<d  <.?:;nI2<d  =.?:;nI2<  >. ?:;nI2<  ?.?:;<cd  @. ?:;n<  A:;  B(   C:;  D:;2  E:;2  F :;I2  G:;2  H.?:;2<d  I I842  J :;I?2<  K :;I?2<  L :;I?2<  M :;I82  N.?:;n2<d  O. ?:;nI2<  P.?:;L2<d  Q :;I?<  R.?:;I<  S.?:;n<  T9:;  U/ I  V.:;I<  W.:;I<  X: :;  Y I  Z. ?:;I<  [I  \!   ]  ^I  _   ` I  a! I/  b.G   c :;I  d  e4 :;I  f :;I  g.G d  h I4  i :;I  j. G   k4 :;I  l.1n@d�B  m 1  n1XY  o�� �B  p.G@�B  q  r4 :;I  s1RUXY  t 1  u 1  vU  w4 1  x.G@d�B  y I4  z :;I  {�� 1  |U  }4 :;I  ~  4 :;I  �4 I  �1RUXY  �1XY  �.G@d�B  � :;I  �4 1  �1RUXY  ��� �B1  �4 :;I  �4 :;I  �4 Gn  �4 G:;n  �.?I4<  �. ?4<  �.?n4<  �.?4<   %U  $ >   :;I  :;   :;I8   I  9:;   :;  	9 :;  
.?:;n<   I  & I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I?<  . ?:;nI<  .?:;nI<d  .?:;n<d   .?:;n<d  !.?:;nI<d  ".?:;nI<d  #.?:;n<  $. ?:;nI<  %.?:;2<d  &.?:;2<cd  '.?:;nI2<d  (.?:;nI2<d  ).?:;n2<d  *.?:;nI2<d  +.?:;nI<  ,/ I  -/ I  . <  /:;  0(   1<  2 :;I?2<  3 :;I?2<  4 :;I?2<  5 :;I2  6:;  7:;2  8.?:;n2<  9:;2  ::;2  ;.?:;nI2<  <.?:;I<  =/ I  ><  ?$ >  @. ?:;I<  A&   B :;n  C9:;  D.?:;n2<d  E :;I82  F.?:;2<cd  G: :;  H I  II  J!   K:;  L! I/  M.G d  N I4  O.G   P :;I  Q :;I  R.G:;@�B  S :;I  T :;I  UU  V4 :;I  W1XY  X 1  Y 1  Z1XY  [ 1  \.G@�B  ]4 :;I  ^4 :;I  _1RUXY  ` 1  a1RUXY  b  c4 :;I  d4 :;I  e4 G:;n  f4 Gn   %U  $ >   :;I  :;   :;I8   I  9:;   :;  	:;  
:;  (   9 :;  .?:;n<   I  & I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d   I8   :;I8  .?:;<d  .?4<d   :;I?2<   :;I?<   . ?:;nI<  !.?:;nI<d  ".?:;n<d  #.?:;n<d  $.?:;nI<d  %.?:;nI<d  &.?:;n<  '. ?:;nI<  (.?:;2<d  ).?:;2<cd  *.?:;nI2<d  +.?:;nI2<d  ,.?:;n2<d  -.?:;nI2<d  ..?:;nI<  // I  0/ I  1 <  2:;  3 :;I?2<  4 :;I?2<  5:;2  6 :;I?<  7.?:;n<d  8:;2  9 I842  : :;I?<  ;. ?:;n<  <.?:;2<cd  =.?:;L2<d  >.?:;n2<  ?.?:;nI2<  @. ?:;nI2<  A:;2  B.?:;<d  C.?:;2<d  D.?:;nI2<d  E. ?:;nI2<  F.?:;<cd  G. ?:;n<  H.?:;I<  I.?:;n<  J.?:;I<  K$ >  L. ?:;I<  M   N:;n  O :;I8  P   Q&   RI  S.?:;I<  T.?:;<  U.?:;<  V :;n  W9:;  X.?:;n2<d  Y/ I  Z:;  [ :;I82  \ :;I2  ]:;  ^.?:;<d  _.?:;nI2<d  `.:;I<  a.:;<  b4 :;I<  c: :;  d I  eI  f!   g:;  h9  i. :;I<  j   k I  l! I/  m.G   n :;I  o  p4 :;I  q.G d  r I4  s4 :;I  t :;I  u :;I  v4 :;I  w4 :;I  x. G   y.G:; d  z :;I  {.1n@d�B  | 1  }���B1  ~�� �B  .G:; d  �1XY  �1XY  � 1  �.G:;@d�B  � I4  �U  �4 :;I  �1XY  � 1  �  �4 1  ��� 1  �1RUXY  � 1  �1RUXY  �1XY  �U  �1RUXY  �1RUXY  �  � 1  �4 1  � :;I  �4 :;I  �.G:;@�B  �.1n@�B  �.G@�B  �. G@�B  �  �.1n@d�B  �4 1  ��� �B1  �.G:;@d�B  � :;I  �4 :;I  �4 :;I  �4 :;I  �.G:;@d�B  � I4  � :;I  ����B  �4 :;I  �4 :;I  �4 G  �4 Gn  �4 G:;n  �4 G:;n  �.?nI4<  �.?n4<  �.?4<  �.?I4<  �. ?4<  �.?4<   %U  $ >   :;I  $ >   I     &   & I  	 :;n  
9:;   :;  9 :;  :;  .?:;n<   I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   :;I8  .?:;2<d   I4  .?:;nI2<d  .?:;n2<d  / I   I82   :;I2  .?:;2<d  :;   I8    :;I8  !.?:;<d  " :;I?2<  # :;I?<  $. ?:;nI<  %.?:;nI<d  &.?:;n<d  '.?:;n<d  (.?:;nI<d  ).?:;nI<d  *.?:;n<  +. ?:;nI<  ,.?:;2<d  -.?:;2<cd  ..?:;nI2<d  /.?:;nI2<d  0.?:;n2<d  1.?:;nI<  2/ I  3 <  4 :;I?2<  5 :;I?2<  6:;2  7 :;I?<  8.?:;<d  9.?:;n<d  ::;2  ;.?:;<d  <.?:;2<d  =.?:;nI2<d  >.?:;nI2<  ?. ?:;nI2<  @.?:;<cd  A. ?:;n<  B:;  C(   D<  E :;I2  F :;I?2<  G :;I?2<  H :;I?2<  I:;  J I842  K :;I82  L.?:;L2<d  M.?:;nLM2<d  N.?:;nILM2<d  O.?:;nILM2<d  P.?:;I<  Q/ I  R9:;  S: :;  T I  U. ?:;I<  VI  W!   XI  Y   Z I  [.G d  \ I4  ].G   ^ :;I  _ :;I  ` :;I  a. G   b  c4 :;I  d :;I  e.1n@d�B  f 1  g1XY  h 1  i 1  j�� �B  k1XY  l��   m�� �B1  n.G@d�B  o I4  p :;I  q :;I  rU  s4 :;I  tU  u4 :;I  v1RUXY  w�� 1  x1XY  y 1  z4 :;I  {.1n@d�B  |4 1  }4 1  ~1XY   1  �4 :;I  � :;I  �4 :;I  �.G@d  � :;I  �4 :;I  �1RUXY  �  �1RUXY  �.1n@d  �.G@d�B  � :;I  ����B  ��� �B  � I4  � :;I  �  � I  �.G@�B  �4 :;I  �4 :;I  �.?I4<  �.?n4<   %U  $ >   :;I  $ >   I     &   & I  	 :;n  
9:;   :;   :;  9 :;  :;  / I  /   /   .?:;n<   I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8    :;I8  !.?:;<d  " :;I?2<  # :;I8  $ :;I?<  %. ?:;nI<  &.?:;nI<d  '.?:;n<d  (.?:;n<d  ).?:;nI<d  *.?:;nI<d  +.?:;n<  ,. ?:;nI<  -.?:;2<d  ..?:;2<cd  /.?:;nI2<d  0.?:;nI2<d  1.?:;n2<d  2.?:;nI2<d  3.?:;nI<  4/ I  5 <  6 :;I?2<  7 :;I?2<  8:;2  9 :;I?<  :.?:;<d  ;.?:;n<d  <:;2  =.?:;<d  >.?:;2<d  ?.?:;nI2<d  @.?:;nI2<  A. ?:;nI2<  B.?:;<cd  C. ?:;n<  D:;  E(   F<  G:;2  H:;2  I :;I2  J:;2  K :;I?2<  L :;I?2<  M :;I?2<  N.?:;n2<d  O:;  P :;I82  Q.?:;n2<d  R.?:;nI2<d  S.?:;2<cd  T.?:;L2<d  U.?:;nILM2<d  V/ I  W.?:;I<  X. ?:;n<  Y9:;  Z.:;<  [.:;<  \: :;  ] I  ^. ?:;I<  _I  `!   a  b.G   c :;I  d.G d  e I4  f :;I  g :;I  h  i4 :;I  j :;I  k4 :;I  l.1n@d�B  m 1  n���B  o�� �B  p1XY  q 1  r��   s�� �B1  t.G@d�B  u I4  v1XY  w :;I  x1XY  y�� 1  z :;I  {���B1  |  }4 1  ~4 :;I  .1n@d�B  �1RUXY  � 1  �1RUXY  �U  �4 1  �.G@d�B  � :;I  � :;I  �.1n@d  �4 :;I  �U  �4 :;I  �1RUXY  �4 1  � 1  �1XY  �4 :;I  �4 :;I  �4 :;I  �. ?4<  �.?n4<   %U  $ >   :;I  :;   :;I8   I  9:;   :;  	9 :;  
.?:;n<   I  & I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I?<  . ?:;nI<  .?:;nI<d  .?:;n<d   .?:;n<d  !.?:;nI<d  ".?:;nI<d  #.?:;n<  $. ?:;nI<  %.?:;2<d  &.?:;2<cd  '.?:;nI2<d  (.?:;nI2<d  ).?:;n2<d  *.?:;nI2<d  +.?:;nI<  ,/ I  -/ I  . <  / :;I?2<  0 :;I?2<  1:;2  2 :;I?<  3.?:;<d  4.?:;n<d  5<  6.?:;2<cd  7.?:;n2<  8. ?:;nI2<  9.?:;nI2<  ::;2  ;.?:;<d  <.?:;2<d  =.?:;nI2<d  >.?:;nI2<  ?.?:;<cd  @. ?:;n<  A:;2  B(   C(   D.?42<d  E:;  F :;I82  G :;I?2<  H :;I2  I.?42<d  J.?:;L2<d  K.?:;nILM2<d  L.?:;nILM2<d  M.?:;I<  N/ I  O.?:;I<  P$ >  Q. ?:;I<  R   S&   T :;n  U9:;  V.?:;n2<d  W:;  X: :;  Y I  ZI  [!   \:;  ].G d  ^ I4  _.4   ` :;I  a :;I  b.G:; d  c.G   d :;I  e.G@d�B  f I4  g I  h :;I  i  j4 :;I  k.1n@d�B  l 1  m1RUXY  n 1  o�� �B  p1XY  q��   r�� 1  s�� �B1  t1RUXY  u4 :;I  v4 :;I  w4 Gn  x.?n4<  y.?:;n<   %U  $ >   :;I  :;   :;I8   I  9:;   :;  	9 :;  
.?:;n<   I  & I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I?<  . ?:;nI<  .?:;nI<d  .?:;n<d   .?:;n<d  !.?:;nI<d  ".?:;nI<d  #.?:;n<  $. ?:;nI<  %.?:;2<d  &.?:;2<cd  '.?:;nI2<d  (.?:;nI2<d  ).?:;n2<d  *.?:;nI2<d  +.?:;nI<  ,/ I  -/ I  . <  / :;I?2<  0 :;I?2<  1:;2  2 :;I?<  3.?:;<d  4.?:;n<d  5<  6.?:;2<cd  7:;2  8.?:;<d  9.?:;2<d  :.?:;nI2<d  ;.?:;nI2<  <. ?:;nI2<  =.?:;<cd  >. ?:;n<  ?:;  @:;2  A:;2  B(   C.?:;nI2<  D<  E0 I  F.?:;n2<d  G.?:;L2<d  H<  I.?:;I<  J$ >  K. ?:;I<  L   M&   N :;n  O9:;  P/ I  Q :;I82  R :;I2  S.?:;2<cd  T: :;  U I  VI  W!   X:;  Y! I/  Z.G d  [ I4  \ :;I  ].G:;@�B  ^ I  _.G@d�B  ` I4  a  b4 :;I  c1XY  d 1  e 1  f1XY  g�� 1  h.1n@d�B  i�� �B  j��   k.1n@d�B  l�� �B1  m4 :;I  n4 :;I  o.?n4<  p.?:;n<   %U  $ >   :;I  ;   $ >   :;I   I     	:;  
 :;I8  I   I  &   & I     :;n  9:;   :;  9:;  :;  .?:;<cd   I4  .?:;n<d  .?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d   <   :;   9 :;  !.?:;n<  ".?:;nI<  #.?:;nI<  $. ?:;nI<  %.?:;nI<  &/ I  ' I82  ( :;I2  ).?:;2<d  *:;  + I8  , :;I8  -.?:;<d  . :;I?2<  / :;I?<  0. ?:;nI<  1.?:;n<d  2.?:;nI<d  3.?:;nI<d  4.?:;n<  5. ?:;nI<  6.?:;2<d  7.?:;2<cd  8.?:;nI2<d  9.?:;nI2<d  :.?:;n2<d  ;/ I  < :;I?2<  = :;I?2<  >:;2  ? :;I?<  @.?:;<d  A.?:;n<d  B:;2  C.?:;<d  D.?:;2<d  E.?:;nI2<d  F.?:;2<cd  G.?:;nI2<  H. ?:;nI2<  I.?:;<cd  J. ?:;n<  K:;  L(   M<  N :;I2  O :;I?2<  P :;I?2<  Q :;I?2<  R.?:;L2<d  S.?:;nILM2<d  T.?:;nILM2<d  U:;2  V(   W.?:;nI2<d  X:;  Y :;I82  Z.?:;nILM2<d  [.?:;nLM2<d  \:;  ].?:;L2<d  ^.?:;n2<d  _.?:;I<  `/ I  a4 :;I<
  b. ?:;n<  c.?:;nI<  d.?:;nI<  e I  fB I  g: :;  h. ?:;I<  iI  j!   k.?:;<  l.?:;I<  m. ?:;I<  n.?:;<  o.G d  p I4  q :;I  r :;I  s.G   t :;I  u. G   v  w4 :;I  x :;I  y4 :;I  z.G@d�B  { I4  | :;I  }1XY  ~ 1  �� 1  �.G@d�B  �U  �4 :;I  �1XY  �1RUXY  �.1n@d�B  � 1  �U  �4 1  �  �4 1  �4 :;I  �1RUXY  �1XY  � 1  �1XY  �1RUXY  ��� �B1  �4 :;I  �4 :;I  �1RUXY  �4 :;I  �  � :;I  �.1n@d�B  ���   � :;I  �4 :;I  �! I/  � 1  � 1  �4 :;I  � I  � I4  �.?4<d  �.?:; d  �.1n@d�B  �4 1  �4 I  ��� �B  ����B1  ��� �B  �4 :;I  �4 :;I  �4 G  �.?I4<  �.?nI4<  �.?n4<  �. ?4<  �.?:;n<   %U  9:;   :;  :;   I8  9 :;   :;   :;I  	.?:;n<  
 I  & I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  9:;  :;   :;I8  .?:;<cd   I4  .?:;n<d  .?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d   <   I82   :;I2  :;2   / I  !:;  " :;I8  #.?:;<d  $.?4<d  %.?4<d  & :;I?2<  ' :;I?<  (. ?:;nI<  ).?:;n<d  *.?:;nI<d  +.?:;nI<d  ,.?:;n<  -. ?:;nI<  ..?:;2<d  /.?:;2<cd  0.?:;nI2<d  1.?:;nI2<d  2.?:;n2<d  3.?:;I<  4.?:;I<  5.?:;nI<  6/ I  7 :;I82  8.?:;2<cd  9.?:;<d  :.?:;nI2<d  ;/ I  < :;I  =4 :;I<
  >   ?.?:;n<  @:;  A :;I82  B :;I2  C.:;I<  D.:;<  E$ >  F$ >  G: :;  H;   I I  J   K&   L :;n  M I  NB I  O. ?:;I<  PI  Q!   R.G   S :;I  T  U4 :;I  V :;I  W.?:;I   X :;I  Y.G d  Z I4  [ :;I  \4 :;I  ]4 :;I  ^.G:; d  _4 :;I  `.G:; d  a. G   b.G:;   c   d  e.1n@d�B  f 1  g1RUXY  h 1  i1RUXY  j1XY  k�� 1  l1XY  mU  n4 1  o.1n@�B  p 1  q�� �B1  r.G@�B  s :;I  t :;I  u :;I  v  w4 1  x. 1n@�B  y.G@d�B  z I4  { :;I  |.G:;@d�B  } I4  ~  4 :;I  �4 :;I  ����B1  ��� �B  �4 :;I  �4 1  �1XY  �1XY  �U  �1RUXY  �.1@d�B  � 1  �1RUXY  � 1  �.G:;@d�B  �4 :;I  � :;I  �4 :;I  ���1  ���   � :;I  � :;I  � I  �4 :;I  �4 :;I  �4 :;I  �4 :;I  �4 G  �4 Gn  �.?I4<  �.?nI4<  �. ?4<  �.?n4<   %U   :;I   I  $ >  ;   $ >      I  	:;n  
 :;I8   :;I8  9:;   :;  9:;  :;  .?:;<cd   I4   I  .?:;n<d  .?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   <   :;  9 :;  :;  .?:;n<   .?:;nI<  !.?:;nI<  ". ?:;nI<  #.?:;nI<  $ I82  % :;I2  &.?:;2<d  ':;  ( I8  ) :;I8  *.?:;<d  +.?4<d  , :;I?2<  - :;I?<  .. ?:;nI<  /.?:;n<d  0.?:;nI<d  1.?:;nI<d  2.?:;n<  3. ?:;nI<  4.?:;2<d  5.?:;2<cd  6.?:;nI2<d  7.?:;nI2<d  8.?:;n2<d  9/ I  :/ I  ;.?:;<d  <.?:;nI2<d  =/ I  > :;I82  ?.?:;nI<cd  @.?:;nI2<cd  A :;  B9 :;  C: :;  Dm:;  E(   F:;  G4 :;I<  H<  I.?42<d  J.?:;I<  K. ?:;n<  L   M.?:;2<d  N.?:;2<cd  O4 :;I<
  P4 :;nI?<  Q4 :;I<
  R   S&   TI  U.?:;I<  V.?:;I<  W.?:;<  X. ?:;I<  Y.?:;<  Z I  [B I  \:;  ] :;I82  ^ :;I2  _.:;I<  `.?:;nI<  a: :;  b :;n  cI  d!   e:;  f.G   g :;I  h  i4 :;I  j.G d  k I4  l4 :;I  m :;I  n.G:; d  o.1@d�B  p 1  q1RUXY  r 1  s1RUXY  tU  u4 1  v�� 1  w.G@�B  x1XY  y :;I  z1RUXY  {1RUXY  |��1  }�� �B  ~ 1  1XY  �1XY  ���   � :;I  �  �4 :;I  �4 :;I  � :;I  �.G@�B  �4 :;I  �4 :;I  �4 G  �4 G  �.?I4<  �.?4<  �  �.?n4<  �.?nI4<   %U  9:;  9:;  :;   :;I8  .?:;<cd   I4   I  	.?:;n<d  
.?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   :;   :;I   <   :;  9 :;  :;  .?:;n<  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<   I82   :;I2  .?:;2<d  :;    I8  ! :;I8  ".?:;<d  #.?4<d  $ :;I?2<  % :;I?<  &. ?:;nI<  '.?:;n<d  (.?:;nI<d  ).?:;nI<d  *.?:;n<  +. ?:;nI<  ,.?:;2<d  -.?:;2<cd  ..?:;nI2<d  /.?:;nI2<d  0.?:;n2<d  1/ I  2/ I  3:;  4(   54 :;I<  6:;  7.?42<d  8.?:;2<cd  9.?:;L2<d  :4 :;I<
  ;   < I  = I  >;   ?B I  @$ >  A$ >  B/ I  C.:;I<  D.:;I<  E: :;  F&   G :;n  H.?:;I<  I. ?:;I<  JI  K!   L.G   M :;I  N  O4 :;I  P.G d  Q I4  R4 :;I  S :;I  T.G:; d  U.1n@d�B  V 1  W���B  X�� �B  Y1XY  Z 1  [��   \�� �B1  ]1RUXY  ^1RUXY  _1XY  `1RUXY  a  b1RUXY  cU  d4 1  e�� 1  f1XY  g 1  h4 1  i4 :;I  j4 :;I  k4 G  l4 G  m.?n4<   %U  9:;  9 :;   :;  :;   :;I  .?:;n<   I  	& I  
.?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;  (   <   :;I2   :;I2   :;I?2<   :;I?2<   :;I?2<  :;2   :;I8  .?:;2<cd   I4  .?:;nI2<d  .?:;nI2<d  / I  / I  .?:;nI2<d  .?:;n2<d   .?:;n2<d  !.?:;n2<d  ".?:;I<  #.?:;I<  $/ I  %9:;  &$ >  '$ >  (: :;  ) :;I  * I  +   , :;I8  -I  .&   /  0 :;n  1 I  2. ?:;I<  3.?:;<  4.?:;I<  5. ?:;I<  6.?:;<  7.G d  8 I4  9 :;I  :.G   ;  <4 :;I  = :;I  >. G   ? :;I  @ :;I  A.G@d�B  B I4  C :;I  DU  E4 :;I  F4 :;I  G4 :;I  H1RUXY  I 1  J  K4 1  L1XY  M  NU  O4 :;I  P4 1  Q1RUXY  R 1  S1RUXY  T1XY  U1XY  V�� 1  W4 I  X��   Y <  Z4 :;I  [4 :;I  \. ?4<  ].?I4<  ^.?n4<   %U  9:;  :;   I82  .?:;2<d   I4  .?:;L2<d  .?:;nILM2<d  	 <  
& I   I  $ >  $ >  .G d   I4  .G@d�B   I4  .1n@d�B   1  ���B  �� �B  1XY   1  ��   �� �B1  .?n4<   I      %U   :;I  $ >  9:;  :;  :;2  (    :;I82  	.?:;nI2<d  
 I4  .?:;nI2<d  <  :;2   :;I8  .?:;<d   I  .?:;<d  .?:;2<d  .?:;nI2<d  & I  .?:;nI2<d  .?:;nILM2<d  :;   I82  .?:;2<cd  .?:;L2<d  .?:;nILM2<d  9  : :;  .:;I<  / I   /   !4 :;I<  " I  # :;  $9:;  %&   &$ >  ' I  (I  )! I/  *.G   + :;I  ,.G d  - I4  .  /4 :;I  04 :;I  1
 :;  2  3 :;I  4 :;I  5 :;I  64 :;I  74 :;I  8.1n@d�B  9 1  :���B  ;�� �B  <1XY  = 1  >��   ?�� �B1  @.1n@d�B  A1RUXY  B�� 1  CU  D4 1  E4 1  F4 1  G1RUXY  H  I1XY  J
 1  KU  L
 1  M  N1XY  O1RUXY  P1XY  Q4 G  R.?n4<  S   T.?nI4<   %U  9 :;  .?:;n@�B   :;I  ���B1  �� �B     .?:;n<  	 I   %U  $ >   :;I  $ >      I  :;n   :;I8  	 :;I8  
9:;   :;   <  .?:;I<   I     & I  &   I  .?:;I<  .?:;I<  .?:;<  . ?:;I<  .?:;<  9:;  :;  4 :;I<   :;  :;n  (     : :;   . G@�B  !4 :;I  "4 :;I  #4 :;I  $4 G   %U  $ >   :;I  $ >      I  :;n   :;I8  	 :;I8  
9:;   :;   <  . ?:;nI<  . ?:;n<  .?:;I<   I     & I  &   I  .?:;I<  .?:;I<  .?:;<  . ?:;I<  .?:;<  :;n  (     :;  9:;  .:;I<   .:;I<  !. ?:;<  "4 :;I<  #. ?:;I<  $ :;  %: :;  &.G   ' :;I  ( :;I  )  *4 :;I  +.G@�B  , :;I  -  .4 :;I  /U  04 :;I  14 :;I  21RUXY  3 1  41XY  54 1  6�� 1  74 :;I  84 :;I  94 G  :.?:;<   %U  $ >  9:;  :;   I842  .?:;L<d   I4  .?:;nLM<d  	:;  
.?:;nLM<d   :;  I     $ >   I   I  9:;  :;   I82  .?:;2<d  .?:;L2<d  .?:;nILM2<d  .?42<d   I  & I   I  .G d   I4  .1n@d�B   1  .G@d�B    I4  !���B1  "�� �B  #.?n4<  $    %U  $ >  9:;   <  & I  <  :;2  (   	9  
: :;  4 :;I<   I   :;  9:;  :;   I842   :;I82  .?:;L2<d   I4  .?:;nI2<d   I  .?:;nILM2<d  .?:;2<cd  .?:;nI<d  .?:;<d  $ >  I      I   I      .G d  ! I4  " :;I  #.1n@d�B  $ 1  %.G@d�B  & I4  ' I  (���B1  )�� �B  * :;I  +1RUXY  , 1  -�� 1  .4 G  /.?n4<  0.?nI4<   %U   :;I  $ >  9:;  :;  :;2  (    :;I82  	.?:;nI2<d  
 I4  .?:;nI2<d  :;  :;2   :;I8  .?:;<d   I  .?:;<d  .?:;2<d  .?:;nI2<d  & I   I82  .?42<d  .?nI42<d  .?:;2<cd  .?:;L2<d  .?:;nILM2<d  .?:;nI2<d  .?:;nILM2<d  <  :;2  9   : :;  !.:;I<  "4 :;I<  # I  $ :;  %9:;  &&   '$ >  ( I  )   *.G d  + I4  , :;I  - :;I  ..G   /.G@d�B  0 I4  1 :;I  2  34 :;I  41XY  5 1  6 1  71RUXY  8 1  9.G@d�B  : I  ;.1n@d�B  <���B  =�� �B  >��   ?�� �B1  @ :;I  A�� 1  B.1n@d  CU  DU  E1XY  F4 G  G.?n4<  H.?nI4<   %U  9:;  :;   I82  .?42<d   I4   I  .?:;2<d  	.?:;L2<d  
.?:;nILM2<d   <  & I   I   I  $ >  $ >  .G d   I4  .G@d�B   I4  .1n@d�B   1  ���B  �� �B  1XY   1  ��   �� �B1  .?:;n<      %U  9:;  9:;  :;   :;I8  .?:;<cd   I4   I  	.?:;n<d  
.?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   :;   :;I   <  . ?:;I<  . ?:;n<  .?:;nI<  .?:;nI<      I   I  ;   B I  $ >  $ >  :;n    :;I8  ! :;I  ":;n  # :;I8  $.?:;I<  %   &&   'I  (.?:;I<  ).?:;I<  *.?:;<  +.?:;<  ,.?:;n<  -4 :;nI?<  .4 :;I<  / :;  0: :;  1.G   2  34 :;I  4.G@�B  5 :;I  6�� 1  7.G@�B  81XY  9  :4 1  ; :;I  <4 :;I  =.1n@�B  >4 1  ?4 :;I  @4 :;I  A4 G  B. ?:;<  C.?I4<  D. ?4<  E.?n4<  F.?4<   %U  $ >  ;   9:;  9:;  :;   :;I8  .?:;<cd  	 I4  
 I  .?:;n<d  .?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   :;   :;I   <  <  .?:;2<d      I   I  B I  $ >  .:;I<  .:;<  . :;<   .?:;I<  !.?:;<  ".?:;<  # :;  $:;  %(   &<  '.?:;2<d  (4 :;I<  ).G d  * I4  +.G   , :;I  -. G   ..G@�B  / :;I  01RUXY  1 1  21XY  31XY  4�� 1  5 :;I  61XY  7 1  8 1  94 G  :.?I4<  ;.?4<  <   %U  $ >   :;I  $ >      I  :;n   :;I8  	 :;I8  
9:;   :;   <  . ?:;n<  .?:;I<   I     & I  &   I  .?:;I<  .?:;I<  .?:;<  . ?:;I<  .?:;<  :;n  (     :;  9:;  4 :;I<   :;   :;  !:;  ".?:;<d  # I4  $.?:;nI<d  %.?:;2<d  &.?:;n2<d  '.?:;nI2<d  ( :;I2  ).?:;2<cd  *.?:;2<d  +4 :;I<  , I  -: :;  .9  /4 :;I<  0.G d  1 I4  2.4   3 :;I  4.G@�B  5 :;I  6
 :;  7U  84 :;I  9  :4 :;I  ;4 :;I  <�� 1  =  >4 :;I  ?�� �B1  @4 :;I  A4 :;I  BI  C! I/  D! I/  E4 G  F4 G  G4 G  H.?:;<   %U  $ >   :;I  ;   $ >      I  :;n  	 :;I8  
 :;I8  9:;   :;  9:;  :;  .?:;<cd   I4   I  .?:;n<d  .?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   <  <  .?:;2<d  . ?:;nI<  .?:;I<      &   !I  ".?:;I<  #.?:;I<  $.?:;<  %. ?:;I<  &.?:;<  ' I  (B I  ).G d  * I4  +.?:;nI@�B  , :;I  -U  .4 :;I  /U  04 :;I  11XY  2 1  3�� 1  44 :;I  54 :;I  6.?I4<  7.?4<  8  9.?:;I<   %U  9:;  :;   I82  .?:;2<d   I4  .?:;L2<d  .?:;nILM2<d  	 <  
& I   I  $ >  $ >  .G d   I4  .G@d�B   I4  .1n@d�B   1  ���B  �� �B  1XY   1  ��   �� �B1  .?n4<   I      %U  $ >  9 :;   :;  9:;  :;   I82  .?:;2<d  	 I4  
.?:;L2<d  9:;   <   I  $ >  .G d   I4  & I  .1n@d�B   1  ���B  �� �B  1XY   1  ��   �� �B1  .?n4<   I      %U  $ >   :;I  9:;  . ?:;<  4 :;I<   :;  $ >  	9:;  
. ?:;n<   I  &   .G@�B  �� 1  4 :;I  & I  4 :;I  4 G  .?:;I<   I   %U   :;I  $ >  9:;  <  :;2  (   :;2  	 :;I8  
.?:;<d   I4   I  .?:;2<d  .?:;nI2<d  & I  9  : :;  :;  .:;I<  /   / I  4 :;I<  .?:;I<   I   :;  9 :;  &   $ >   I  .G    :;I   .G d  ! I4  "   #.G@�B  $ :;I  %U  &4 :;I  '4 :;I  (4 :;I  )1RUXY  * 1  + 1  ,1XY  -1RUXY  . 1  /  04 G   %U  9:;  9:;  :;   :;I8  .?:;<cd   I4   I  	.?:;n<d  
.?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   :;   :;I   <  <  .?:;2<d  <      I   I  ;   B I  $ >  $ >  :;n   :;I8    :;I  !:;n  " :;I8  #.?:;I<  $   %&   &I  '.?:;I<  (.?:;I<  ).?:;<  *. ?:;I<  +.?:;<  ,. ?:;<  -4 :;I<  . :;  /  0.G d  1 I4  2.G@�B  31XY  4 1  5�� 1  64 :;I  74 :;I  84 G  9.?I4<  :.?4<   %U   :;I  $ >  9:;  <  :;2  (   :;2  	 :;I8  
.?:;<d   I4   I  .?:;<d  .?:;2<d  .?:;nI2<d  & I  .?:;nILM2<d  :;2  9  : :;  .:;I<  /   4 :;I<  :;   I82   :;I82  .?:;2<cd  .?:;L2<d  .?:;2<d  .?:;nI2<d  .?:;nILM2<d   .?:;nILM2<d  ! I  " :;  #9:;  $&   %$ >  & I  '.G d  ( I4  ) :;I  *.G   + :;I  ,.1n@d�B  - 1  .���B  /�� �B  01XY  1 1  2��   3�� �B1  4.G@d  5 I4  6 :;I  7�� 1  81XY  9.1n@d  :U  ;4 G  <.?n4<  =   >.?nI4<   %  $ >  $ >   :;I  9:;  4 :;nI?<  4 :;I<   :;  	9:;  
 I     4 G  & I  4 G   %U  $ >   :;I  $ >      :;I   I  :;n  	 :;I8  
 :;I8  9:;   :;  <  .?:;nI2<d   I4  & I   <  .?:;I<   I     &   I  .?:;I<  .?:;I<  .?:;<  . ?:;I<  .?:;<  9:;  . ?:;I<   :;  :;     !: :;  ".G d  # I4  $. ?:;n<  %.G@�B  &  '4 :;I  (4 :;I  )U  *4 :;I  +1RUXY  , 1  -�� 1  . I  /4 :;I  04 :;I  14 :;I?<  2.?nI4<  3.?I4<  4. ?4<  5. ?:;<  6.?n4<   %U  $ >  9:;  :;   :;I8  .:;I<   I  .:;I<  	. ?:;I<  
4 :;I<  . ?:;I<   :;   :;I  $ >  :;n  (    I       9:;   <     & I  .G    :;I   :;I  .G@�B  U  4 :;I    4 :;I   1XY  ! 1  "�� 1  #4 G   %  $ >  $ >   :;I  9:;  4 :;nI?<  4 :;I<   :;  	9:;  
 I     4 G  & I  4 G   %U  9:;  9:;  :;   :;I8  .?:;<cd   I4   I  	.?:;n<d  
.?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   :;   :;I   <  :;   I82  .?:;L2<d  .?:;nILM2<d      I   I  ;   B I  $ >  $ >  .G d    I4  !.G@d�B  " I4  #.1n@d�B  $ 1  %���B  &�� �B  '1XY  ( 1  )��   *�� �B1  +.?:;n<   %U  $ >   :;I  :;   :;I8   I  9:;   :;  	9 :;  
.?:;n<   I  & I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d  .?4<d   :;I?2<   :;I?<  . ?:;nI<  .?:;nI<d   .?:;n<d  !.?:;n<d  ".?:;nI<d  #.?:;nI<d  $.?:;n<  %. ?:;nI<  &.?:;2<d  '.?:;2<cd  (.?:;nI2<d  ).?:;nI2<d  *.?:;n2<d  +.?:;nI2<d  ,.?:;nI<  -/ I  ./ I  / <  0 :;I?2<  1 :;I?2<  2:;2  3 :;I?<  4.?:;<d  5<  6.?:;2<cd  7. ?:;nI2<  8:;2  9.?:;<d  :.?:;2<d  ;.?:;nI2<d  <.?:;nI2<  =.?:;<cd  >. ?:;n<  ?.?42<d  @:;  A:;2  B :;I?2<  C<  D :;I2  E.?:;n2<d  F0 I  G.?:;I<  H.?:;<d  I.?:;I<  J$ >  K. ?:;I<  L   M:;n  N :;I8  O   P&   QI  R.?:;I<  S.?:;<  T.?:;<  U :;n  V9:;  W.?:;n2<d  X/ I  Y :;I82  Z:;  [(   \.?:;nI2<d  ].:;I<  ^.:;<  _4 :;I<  `: :;  a I  bI  c!   d:;  e! I/  f9  g. :;I<  h4 :;I<  i.G   j :;I  k  l4 :;I  m.G d  n I4  o4 :;I  p :;I  q.?:;I   r.?:;   s :;I  t.G:; d  u.G:; d  v. G:;   w.1@�B  x  y4 1  z�� 1  { :;I  |4 :;I  }  ~4 :;I  .1n@d�B  � 1  �U  �4 1  �  �1XY  � 1  �1RUXY  ���   �1XY  �1XY  �.1n@�B  ��� �B1  �1RUXY  �.G:;@�B  �.G:;@�B  � :;I  �4 :;I  �4 :;I  �1XY  �1RUXY  �1RUXY  �U  � 1  �4 1  �4 :;I  �4 :;I  �4 G  �! I/  �4 G  �4 G:;n  �.?I4<  �.?4<  �.?n4<  �.?4<   %U  $ >   :;I  $ >   I     &   & I  	 :;n  
9:;   :;  9 :;  :;  .?:;n<   I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d  .?4<d   :;I?2<    :;I8  ! :;I?<  ". ?:;nI<  #.?:;nI<d  $.?:;n<d  %.?:;n<d  &.?:;nI<d  '.?:;nI<d  (.?:;n<  ). ?:;nI<  *.?:;2<d  +.?:;2<cd  ,.?:;nI2<d  -.?:;nI2<d  ..?:;n2<d  /.?:;nI2<d  0.?:;nI<  1/ I  2/ I  3 <  4:;  5(   6<  7:;2  8.?42<d  9.?:;L2<d  :.?:;nILM2<d  ; :;I?2<  < :;I?2<  = :;I?2<  > :;I2  ?9:;  @.?:;n2<d  A/ I  B.:;I<  C.:;I<  D: :;  E I  F.?:;I<  G. ?:;I<  HI  I!   J.G   K :;I  L  M4 :;I  N.G d  O I4  P4 :;I  Q :;I  R.G:; d  S.G@d�B  T I4  U.1n@d�B  V 1  W1RUXY  X 1  Y1RUXY  Z1XY  [1RUXY  \  ] 1  ^1RUXY  _U  `4 1  a�� 1  b��   c�� �B1  d4 :;I  e4 :;I  f.?n4<  g.?4<   %U  $ >   :;I  :;   :;I8   I  9:;   :;  	9 :;  
.?:;n<   I  & I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I?<  . ?:;nI<  .?:;nI<d  .?:;n<d   .?:;n<d  !.?:;nI<d  ".?:;nI<d  #.?:;n<  $. ?:;nI<  %.?:;2<d  &.?:;2<cd  '.?:;nI2<d  (.?:;nI2<d  ).?:;n2<d  *.?:;nI2<d  +.?:;nI<  ,/ I  -/ I  . <  / :;I?2<  0 :;I?2<  1:;2  2 :;I?<  3.?:;<d  4.?:;n<d  5<  6.?:;2<cd  7:;2  8.?:;<d  9.?:;2<d  :.?:;nI2<d  ;.?:;nI2<  <. ?:;nI2<  =.?:;<cd  >. ?:;n<  ? :;I?<  @ :;I?<  A.?4<d  B. ?:;nI2<  C.?:;nILM2<d  D.?:;nILM2<d  E.?:;I<  F$ >  G. ?:;I<  H   I&   J :;n  K9:;  L.?:;n2<d  M/ I  N:;  O :;I82  P :;I2  Q.?:;2<cd  R: :;  S I  TI  U!   V:;  W:;n  X :;I8  Y   ZI  [.?:;I<  \.?:;I<  ].?:;<  ^.?:;<  _.G d  ` I4  a :;I  b.G:; d  c. G   d. 1n@�B  e :;I  f.1n@d�B  g 1  h 1  i1RUXY  j.G@d�B  k I4  l :;I  m�� 1  n :;I  o :;I  p4 :;I  q4 :;I  r.?:;I<   %U  $ >   :;I  :;   :;I8   I  9:;   :;  	9 :;  
<  .?:;nI2<d   I4   I  / I  & I  .?:;I<  $ >  . ?:;I<   :;n  9:;  : :;  :;  .G@d�B   I4   :;I  U  4 :;I  �� 1   I4   :;I   :;I   ���B1  !�� �B  "4 :;I  #4 :;I   %  $ >   :;I  $ >   :;I   I     :;  	 :;I8  
I   I  &   & I     :;n  9:;   :;  9 :;  4 :;nI?<  4 :;nI?<  9:;  : :;  .?:;I<  . ?:;I<  .?:;<  .?:;I<  . ?:;I<  .?:;<  4 :;I  4 :;I  I   ! I/  !4 G   %U  $ >   :;I  $ >   I     &   & I  	 :;n  
9:;   :;  9 :;  :;  .?:;n<   I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  <  .?:;L2<d   I4  .?:;2<cd   :;I2  .?:;2<d  / I  / I  :;   :;I82  :;   I82   .?:;2<cd  !.?:;L2<d  ".?:;n2<d  #.?:;nI<  $ :;I8  %.?:;I<  &. ?:;I<  '9:;  (: :;  ) I  *.G d  + I4  , :;I  -.1n@d�B  . 1  /1XY  0�� �B  1 1  21XY  3��   4�� �B1  5.G@�B  6 :;I  7 :;I  8�� 1  91RUXY  : 1  ;4 :;I  <4 :;I  =.?n4<   %U  $ >   :;I  :;   :;I8   I  9:;   :;  	9 :;  
.?:;n<   I  & I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I?<  . ?:;nI<  .?:;nI<d  .?:;n<d   .?:;n<d  !.?:;nI<d  ".?:;nI<d  #.?:;n<  $. ?:;nI<  %.?:;2<d  &.?:;2<cd  '.?:;nI2<d  (.?:;nI2<d  ).?:;n2<d  *.?:;nI2<d  +.?:;nI<  ,/ I  -/ I  . <  / :;I?2<  0 :;I?2<  1:;2  2 :;I?<  3.?:;<d  4.?:;n<d  5<  6.?:;2<cd  7:;2  8.?:;<d  9.?:;2<d  :.?:;nI2<d  ;.?:;nI2<  <. ?:;nI2<  =.?:;<cd  >. ?:;n<  ?<  @.?:;n2<d  A.?:;L2<d  B.?:;I<  C$ >  D. ?:;I<  E   F&   G :;n  H9:;  I/ I  J:;  K :;I82  L :;I2  M.?:;2<cd  N: :;  O I  PI  Q!   R:;  S.G d  T I4  U :;I  V.G@d�B  W I4  X I  Y  Z4 :;I  [1XY  \ 1  ] 1  ^1XY  _�� 1  `.1n@d�B  a�� �B  b��   c.1n@d�B  d�� �B1  e4 :;I  f4 :;I  g.?n4<  h.?:;n<   %U  $ >   :;I  $ >   I     &   & I  	 :;n  
9:;   :;   :;  9 :;  :;  .?:;n<   I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   :;I8  .?:;2<d   I4  .?:;nI2<d  .?:;n2<d  / I   I82   :;I2  .?:;2<d  :;    I8  ! :;I8  ".?:;<d  #.?4<d  $ :;I?2<  % :;I?<  &. ?:;nI<  '.?:;nI<d  (.?:;n<d  ).?:;n<d  *.?:;nI<d  +.?:;nI<d  ,.?:;n<  -. ?:;nI<  ..?:;2<d  /.?:;2<cd  0.?:;nI2<d  1.?:;nI2<d  2.?:;n2<d  3.?:;nI<  4/ I  5 <  6 :;I?2<  7 :;I?2<  8:;2  9 :;I?<  :.?:;n<d  ;<  <.?:;2<cd  =:;2  >.?:;<d  ?.?:;2<d  @.?:;nI2<d  A.?:;nI2<  B. ?:;nI2<  C.?:;<cd  D. ?:;n<  E:;  F(   G :;I2  H :;I?2<  I :;I?2<  J :;I?2<  K :;I?<  L :;I?<  M.?:;nI2<d  N:;  O I8L2  P I842  Q :;I82  R.?:;L2<d  S.?:;nI2<d  T.?:;nILM2<d  U.?:;L2<d  V.?:;n2<d  W.?4<d  X/ I  Y<  Z.?:;I<  [ :;I?2<  \. ?:;n<  ]9:;  ^.:;I<  _.:;I<  `: :;  a I  b. ?:;I<  cI  d!   eI  f   g I  h.G   i :;I  j  k4 :;I  l.G d  m I4  n4 :;I  o :;I  p4 :;I  q :;I  r :;I  s. G   t.G:; d  u.G:; d  v.1n@d�B  w 1  x 1  y1XY  z�� �B  {1XY  |1RUXY  }��   ~�� �B1  ���B1  ��� �B  ��� 1  �.G@d�B  � I4  � :;I  ����B�B  �.G@d�B  � :;I  �1RUXY  � 1  �1RUXY  �  �1XY  �.1n@d�B  �U  �4 1  �U  �4 1  �1RUXY  �1XY  � 1  �  �.G:;@d�B  � :;I  �4 :;I  �4 :;I  �4 :;I  �4 I  �.G:;@d�B  � :;I  �4 :;I  �4 :;I  �.G:;@d�B  �4 :;I  �4 :;I  � :;I  �4 :;I  �4 :;I  � 1  �4 :;I  �.G@�B  � :;I  �.G@�B  � :;I  � :;I  �4 :;I  �.?n4<  �. ?4<  �.?I4<   %U  $ >   :;I  $ >   I  &   & I   :;n  	9:;  
 :;  9 :;  :;  .?:;n<   I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I8   :;I?<   . ?:;nI<  !.?:;nI<d  ".?:;n<d  #.?:;n<d  $.?:;nI<d  %.?:;nI<d  &.?:;n<  '. ?:;nI<  (.?:;2<d  ).?:;2<cd  *.?:;nI2<d  +.?:;nI2<d  ,.?:;n2<d  -.?:;nI2<d  ..?:;nI<  // I  0/ I  1 <  2 :;I?2<  3 :;I?2<  4:;2  5 :;I?<  6.?:;<d  7.?:;n<d  8:;2  9.?:;<d  :.?:;2<d  ;.?:;nI2<d  <.?:;nI2<  =. ?:;nI2<  >.?:;<cd  ?. ?:;n<  @:;  A(   B<  C:;2  D.?:;n2<d  E :;I?2<  F :;I?2<  G :;I?2<  H :;I2  I.?:;n2<d  J.?:;I<  K9:;  L/ I  M:;  N :;I82  O.?:;2<cd  P: :;  Q I  R.?:;I<  S. ?:;I<  TI  U!   V:;  W.G   X :;I  Y.G@d�B  Z I4  [��   \�� 1  ] :;I  ^  _4 :;I  `4 :;I  a4 :;I   %U  $ >   :;I  $ >      :;I   I  :;  	 :;I8  
I   I  &   & I    9:;   :;  9 :;  :;  (   <   :;I2   :;I2   :;I?2<   :;I?2<   :;I?2<  :;  .?:;2<d   I4  .?:;nI2<d  .?:;nI2<d  .?:;nI2<d   :;  ! :;I?<  ". ?:;nI<  #. ?:;nI<  $.?:;<  %.?:;I<  &.?:;I<  '. ?:;I<  (.?:;<  ). ?:;I<  * :;n  +9:;  ,: :;  -9  ..:;I<  /.:;I<  0.G   1 :;I  2   3.G:; d  4 I4  5. G   6.G:; d  7.G@�B  8 :;I  9 :;I  :U  ;4 :;I  <�� 1  =.1n@d�B  > 1  ?.G:;@d�B  @ I4  A :;I  B I  C  D1XY  E 1  FU  G4 :;I  H1RUXY  I U  J.G:;@d�B  K4 :;I  L1XY  M���B1  N�� �B  O :;I  P :;I  Q��1  R��1  S�� �B1  T4 :;I  U4 :;I  V4 :;I  W4 :;I?<  X.?n4<  Y.?4<   %U  $ >   :;I  :;   :;I8   I  9:;   :;  	9 :;  
.?:;n<   I  & I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I?<  . ?:;nI<  .?:;nI<d  .?:;n<d   .?:;n<d  !.?:;nI<d  ".?:;nI<d  #.?:;n<  $. ?:;nI<  %.?:;2<d  &.?:;2<cd  '.?:;nI2<d  (.?:;nI2<d  ).?:;n2<d  *.?:;nI2<d  +.?:;nI<  ,/ I  -/ I  . <  / :;I  0<  1.?:;nILM2<d  2.?:;I<  3$ >  4. ?:;I<  5&   6 :;n  79:;  8.?:;n2<d  9/ I  ::;  ; :;I82  < :;I2  =.?:;2<cd  >: :;  ? I  @I  A!   B:;  C.G@d�B  D I4  E I  F :;I  G��   H4 :;I  I4 :;I   %U  9:;  9 :;   :;  :;   :;I  .?:;n<   I  	& I  
.?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d  .?4<d   :;I?2<   :;I8   :;I?<  . ?:;nI<  .?:;nI<d  .?:;n<d  .?:;n<d   .?:;nI<d  !.?:;nI<d  ".?:;n<  #. ?:;nI<  $.?:;2<d  %.?:;2<cd  &.?:;nI2<d  '.?:;nI2<d  (.?:;n2<d  ).?:;nI2<d  *.?:;nI<  +/ I  ,/ I  - <  .:;  /.?42<d  0.?:;L2<d  1.?:;L2<d  2.?:;nILM2<d  3<  49:;  5.?:;n2<d  6/ I  7.:;I<  8.:;I<  9$ >  :$ >  ;: :;  < I  =   >&   ? :;n  @ I  A.?:;I<  B. ?:;I<  CI  D!   E.G   F :;I  G  H4 :;I  I.G d  J I4  K4 :;I  L :;I  M.G:; d  N.G@d�B  O I4  P.1n@d�B  Q 1  R1RUXY  S 1  T1RUXY  U1XY  V1RUXY  W  X 1  Y1RUXY  ZU  [4 1  \�� 1  ]��   ^���B1  _�� �B  `1XY  a�� �B1  b4 :;I  c4 :;I  d.?n4<   %U  9:;   :;  9 :;  :;   :;I  .?:;n<   I  	& I  
.?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I8   :;I?<  . ?:;nI<  .?:;nI<d  .?:;n<d  .?:;n<d  .?:;nI<d   .?:;nI<d  !.?:;n<  ". ?:;nI<  #.?:;2<d  $.?:;2<cd  %.?:;nI2<d  &.?:;nI2<d  '.?:;n2<d  (.?:;nI2<d  ).?:;nI<  */ I  +/ I  , <  - :;I?2<  . :;I?2<  /:;2  0 :;I?<  1.?:;<d  2.?:;n<d  3<  4.?:;n2<  5.?:;nI2<  6.?:;nI2<  7:;2  8.?:;<d  9.?:;2<d  :.?:;nI2<d  ;.?:;nI2<  <. ?:;nI2<  =.?:;<cd  >. ?:;n<  ?:;  @(   A :;I2  B :;I?2<  C :;I?2<  D :;I?2<  E :;I?<  F :;I?<  G :;I?<  H.?:;n<  I9:;  J.?:;n2<d  K/ I  L:;  M :;I82  N.?:;2<cd  O4 :;I<  P$ >  Q$ >  R   S :;I  T I  U:;n  V :;I8  W.?:;I<  X   Y&   ZI  [.?:;I<  \.?:;I<  ].?:;<  ^. ?:;I<  _.?:;<  `  a. ?:;I<  b :;n  c: :;  d I  eI  f!   g:;  h. G   i.G@�B  j :;I  k :;I  l I  mU  n4 :;I  o4 :;I  p�� 1  q4 :;I  r�� �B1  s :;I  t4 :;I  u4 :;I  v! I/  w4 G  x4 G:;n  y.?I4<  z.?n4<  {.?4<  |.?:;I<  }    %U  $ >   :;I  :;   :;I8   I  9:;   :;  	9 :;  
.?:;n<   I  & I  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<  :;   I82   :;I2  .?:;2<d   I4  .?:;2<d  :;   I8   :;I8  .?:;<d   :;I?2<   :;I?<  . ?:;nI<  .?:;nI<d  .?:;n<d   .?:;n<d  !.?:;nI<d  ".?:;nI<d  #.?:;n<  $. ?:;nI<  %.?:;2<d  &.?:;2<cd  '.?:;nI2<d  (.?:;nI2<d  ).?:;n2<d  *.?:;nI2<d  +.?:;nI<  ,/ I  -/ I  . <  / :;I?2<  0 :;I?2<  1:;2  2 :;I?<  3.?:;<d  4.?:;n<d  5<  6.?:;2<cd  7:;2  8.?:;<d  9.?:;2<d  :.?:;nI2<d  ;.?:;nI2<  <. ?:;nI2<  =.?:;<cd  >. ?:;n<  ?.?:;n2<d  @<  A.?:;<d  B.?:;I<  C$ >  D. ?:;I<  E   F&   G :;n  H9:;  I/ I  J:;  K :;I82  L :;I2  M.?:;2<cd  N: :;  O I  PI  Q!   R:;  S:;n  T :;I8  U   VI  W.?:;I<  X.?:;I<  Y.?:;<  Z.?:;<  [.G d  \ I4  ] :;I  ^.G@d�B  _ I4  ` :;I  a :;I  b  c4 :;I  d�� 1  e :;I  f I  g1XY  h 1  i 1  j1XY  k4 :;I  l4 :;I  m.?I4<  n.?n4<  o.?4<  p.?:;nI<   %U  9:;  9:;  :;   :;I8  .?:;<cd   I4   I  	.?:;n<d  
.?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   :;   :;I   <   :;  9 :;   :;  :;   I82  .?42<d  .?:;L2<d  .?:;nILM2<d  4 :;I<
  4 :;I<
      I    I  !;   "B I  #$ >  $$ >  %: :;  & :;n  ':;  (.?:;I<  ). ?:;I<  *.G d  + I4  ,.G@d�B  - I4  ..1n@d�B  / 1  0���B  1�� �B  21XY  3 1  4��   5�� �B1  64 :;I  74 :;I  84 G  9.?:;n<   %U  $ >   :;I   I  9:;   :;   :;  9 :;  	9:;  
:;   :;I8  .?:;<cd   I4   I  .?:;n<d  .?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   <  :;  (   <   :;I2   :;I?2<   :;I?2<   :;I?2<   :;I2   .?:;I<  !4 :;I<
  ".?:;n<  #.?:;nI<  $/ I  %$ >  &;   ' I  (   )&   * :;n  +:;  ,. ?:;I<  -.?:;nI<  ..?:;nI<  /: :;  0 I  1B I  2.G   3 :;I  4.G@�B  5 :;I  6U  74 :;I  84 :;I  94 :;I  :4 :;I  ;�� 1  <I  =! I/  > :;I  ?4 :;I  @U  A  B4 :;I  C4 G  D.?I4<   %U  9:;  9:;  :;   :;I8  .?:;<cd   I4   I  	.?:;n<d  
.?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   :;   :;I   <   :;  9 :;  :;  .?:;n<  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<   I82   :;I2  .?:;2<d  :;    I8  ! :;I8  ".?:;<d  #.?4<d  $ :;I?2<  % :;I?<  &. ?:;nI<  '.?:;n<d  (.?:;nI<d  ).?:;nI<d  *.?:;n<  +. ?:;nI<  ,.?:;2<d  -.?:;2<cd  ..?:;nI2<d  /.?:;nI2<d  0.?:;n2<d  1/ I  2/ I  3.?:;<d  4.?:;nI2<d  5/ I  6 :;  79 :;  8: :;  9 :;I82  :.?:;nI<cd  ;.?:;nI2<cd  <:;  =(   >m:;  ?:;  @.?:;2<cd  A.?:;L2<d  B.?:;nILM2<d  C4 :;nI?<  D4 :;I<
  E4 :;I<
  F   G I  H I  I;   JB I  K$ >  L$ >  M:;  N :;I82  O :;I2  P4 :;I<  Q.:;I<  R.:;I<  S: :;  T&   U :;n  V.?:;I<  W. ?:;I<  XI  Y!   Z:;  [9  \:;  ].4<d  ^.:;ILM<d  _.L4<d  `. :;I<  a.G   b :;I  c  d4 :;I  e.G d  f I4  g4 :;I  h.G:; d  i :;I  j :;I  k.G:; d  l :;I  m. G   n.G@d�B  o I4  p.1@d�B  q 1  r���B  s�� �B  t1XY  u 1  v��   w�� �B1  x.1n@d�B  y 1  z.G@d�B  {1RUXY  |1RUXY  }U  ~4 1  1XY  ��� 1  �1RUXY  �  �1XY  � 1  �4 1  �1RUXY  �4 1  �U  �.G@�B  �4 :;I  �4 :;I  �4 I?4<  �4 G  �4 G  �.?n4<  �.?I4<  �.?4<  �   %U  $ >   :;I  ;   9:;   :;  9:;  :;  	 :;I8  
.?:;<cd   I4   I  .?:;n<d  .?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   <   :;  9 :;  :;  .?:;n<  .?:;nI<  .?:;nI<  . ?:;nI<  .?:;nI<   I82   :;I2   .?:;2<d  !:;  " I8  # :;I8  $.?:;<d  % :;I?2<  & :;I?<  '. ?:;nI<  (.?:;n<d  ).?:;nI<d  *.?:;nI<d  +.?:;n<  ,. ?:;nI<  -.?:;2<d  ..?:;2<cd  /.?:;nI2<d  0.?:;nI2<d  1.?:;n2<d  2/ I  3/ I  4.?:;<d  5.?:;nI2<d  6/ I  7:;  8 I842  9.?:;L2<d  :.?:;nILM2<d  ; :;I82  <.?:;nI<cd  =.?:;nI2<cd  >:;  ?.?:;L2<d  @.?:;nI2<d  A.?:;I<  B4 :;I<
  C.?:;I<  D$ >  E I  F   G&   H :;n  I I  JB I  K:;  L :;I82  M :;I2  N: :;  O. ?:;I<  PI  Q!   R9  S:;  T.4<d  U.:;ILM<d  V.L4<d  W4 :;I<  XI  Y   Z I  [.G d  \ I4  ] :;I  ^ :;I  _.G   ` :;I  a.G:; d  b.4   c.G@d�B  d I4  e.1n@d�B  f 1  g1XY  h :;I  i :;I  j.1@d�B  k���B1  l�� �B  m�� 1  n��   o���B  p1XY  q 1  r�� �B1  s.G@d�B  t1XY  u 1  v1RUXY  w. G@�B  x.G:;@d�B  y.4@�B  z 1  { 1  |4 :;I  }4 :;I  ~4 I?4<  4 G  �4 G  �.?I4<  �   %U  9:;  9:;  :;   :;I8  .?:;<cd   I4   I  	.?:;n<d  
.?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   :;   :;I   <   :;  .?:;nI<  . ?:;nI<  4 :;nI?<
      I   I  ;   B I  $ >  $ >      9  !4 :;I<  ": :;  #.G@�B  $ :;I  %  &4 :;I  '4 G   %U  9:;  9:;  :;   :;I8  .?:;<cd   I4   I  	.?:;n<d  
.?:;nI<d  .?:;2<d  .?:;nI2<d  .?:;n2<d  .?:;nI2<cd  .?:;nI2<d  & I   :;   :;I   <  :;   I82  .?:;L2<d  .?:;nILM2<d      I   I  ;   B I  $ >  $ >  .G d    I4  !.G@d�B  " I4  #.1n@d�B  $ 1  %���B  &�� �B  '1XY  ( 1  )��   *�� �B1  +.?:;n<   %  $ >   :;I  $ >      I  &   & I  	'  
 I  :;  (   :;   :;I8  :;   :;I8   :;I8   :;I8  :;  :;   :;I  :;  :;   :;I8   :;I8  I  ! I/  .:;'I    :;I  4 :;I   :;I   4 :;I  !.:;'   "  #! I  $.:;'I@�B  % :;I  & :;I  '1RUXY  ( 1  )U  *4 1  + :;I  ,1XY  -  .1XY  /.:;'I@�B  04 :;I  14 :;I  24 :;I  34 :;I  4��1  5�� �B  6 :;I  7U  8  91RUXY  :4 1  ;.:;'@�B  <
 :;  =.1@�B  >.1@�B  ? 1  @�� 1�B  A�� 1  B 1  C��1  D4 1  E.:;'@�B  F�� �B1  G���B1  H  I 1  J4 1I  K4 4I  L! I/  M.?:;'I@�B  N4 :;I  O4 :;I  P.?:;'I<  Q.?:;'<  R.?'I4<  S.?:;'I<  T   U.?:;'I<   %  $ >  $ >   :;I  :;   :;I8   :;I8  :;  	 :;I  
 :;I  .:;'I    :;I  4 :;I     I  & I  .?:;'I@�B   :;I  1RUXY   1   1   1  U  4 1  4 1  4 :;I  4 :;I   %  $ >  $ >   :;I  :;   :;I8   :;I8  :;  	 :;I  
 :;I  .:;'I    :;I  4 :;I     I  & I  .?:;'I@�B   :;I  4 :;I  1RUXY   1   1  U  4 1  4 1    4 :;I  4 :;I   %  $ >   :;I  $ >      I  &   & I  	:;  
(   :;  '   I  :;   :;I8  'I   :;I8   :;I  I  ! I   :;I  :;   :;I   :;I  :;  ! I/  :;  :;   :;I8   :;I8  :;    :;I  ! :;I  ".:;'I   # :;I  $.:;'   % :;I  &4 :;I  '.:;'   ( :;I  ) :;I  *.:;'I   +.?:;'I   ,4 :;I  -. :;'   ..:;'I@�B  / :;I  04 :;I  1  2  3.:;'@�B  4 :;I  5 :;I  64 :;I  71RUXY  8 1  9U  :4 :;I  ;4 :;I  <4 1  =U  >4 :;I  ?1RUXY  @1XY  A1XY  B  C4 1  D 1  E  F4 1  G��1  H�� �B  I1XY  J1XY  K�� 1  L��1  M4 :;I  N.:;'I@�B  O.?:;'I   P :;I  Q
 :;  R 1  S 1  T1RUXY  U4 :;I  V 1XY  W.:;'I@�B  X :;I  Y4 :;I  Z�� �B  [.1@�B  \.?:;'@�B  ] :;I  ^.?:;'I@�B  _.?:;'I@�B  `4 :;I  a1RUXY  b.?:;'I@�B  c.?:;'@�B  d.?:;'@�B  e.?:;'I@�B  f4 :;I  g4 :;I  h. ?:;'<  i.?:;'I<   %  $ >   :;I  $ >      I  &   & I  	:;  
(    :;I  :;   :;I8  I  ! I  :;   :;I  :;   :;I8   :;I   :;I8   :;I  'I   I  :;   :;I8  .:;'I    :;I   :;I  .:;'I    :;I   .:;'   ! :;I  "4 :;I  #  $4 :;I  %4 :;I  &.?:;'   '.?:;'I   (.:;'I@�B  ) :;I  *4 :;I  +.:;'I@�B  , :;I  -4 :;I  ..:;'@�B  / :;I  0 :;I  14 :;I  2U  3�� �B  4 :;I  5��1  6�� �B  7��1  8 :;I  9�� 1  : :;I  ;:;  <4 :;I  =  >4 :;I  ?1XY  @ 1  A 1  B  C4 1  D4 :;I  E4 :;I  F1XY  G4 1  H1RUXY  I1XY  J.:;'I@�B  K4 :;I  L
 :;  M  NU  O4 1  P
 1  Q1RUXY  R.1@�B  S1XY  T 1  U.?:;'@�B  V :;I  W1RUXY  X 1  Y.?:;'I@�B  Z
 :;  [���B1  \.?:;'I@�B  ]4 :;I  ^4 :;I  _4 :;I  `. ?:;'<  a.?:;'I<  b.?:;'<   �   �  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include  del_op.cc   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   cstdlib   <built-in>    malloc.h     ��, �   ?  �      /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/../libgcc ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include  unwind-pe.h   eh_personality.cc   unwind-cxx.h   exception   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   cstdlib   cxxabi.h   unwind.h   <built-in>      ��]* � u u ; +	J XY�0  0���lɠLk  ����q.J	f)�/<LYu-/K2hm�/=v�==k��I1k���uu;+� �==�H�� <�J=/� <0
  ��� MkJ[�wi��r�   ���IK��*�uu;+� JNz ��t<.  ��� =M
J�v�
.q����yJ�  �2j*\*N . � M 9 1 K���~��<�~<�-=� fuu;+@J�8�*L.; uu;+IJ�h��   ��=.CX<XDX��+��.�}J� f�X� f�� �u� ����!�v!%Y�}Ȇ
 1�Y:L83#��~��~a�.�~��uu;+�JR�>.� X8J��^zX�}fvI>G>A8��ts�Z�x.ut�~ r��tfX�~��K-/gJs.f4�L��Z��~.��Lyt Xn��I/Z�.KIYu �}� �~f *�uu;+�J �XJ�	<OXy� J��"�K�����>J��F��~�.$��   ���@f==:?i��Y�}.���wqtnX(���z��f�	 �    �   �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits  new_opv.cc   <built-in>    c++config.h   new     �g��	 �     �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include  eh_throw.cc   unwind-cxx.h   exception_ptr.h   cstddef   c++config.h   exception   stddef.h   unwind.h   atomic_word.h   <built-in>    cxxabi.h      � 	JwX	J2w=;K�NF�sX  p�=JMYPItv<=u�YeCz<uyj�  ��� KY0M�J�~ Yf��iX\    �  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  eh_call.cc   unwind-cxx.h   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   cstdlib   exception   unwind.h   cxxabi.h   <built-in>      @�'JLM���}���    A  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext  locale_facets.h   ostream   basic_ios.h   streambuf   ios_base.h   ostream.tcc   postypes.h   streambuf.tcc   char_traits.h   iomanip   ostream_insert.h   streambuf_iterator.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   stl_iterator_base_types.h   c++config.h   cwchar   clocale   allocator.h   basic_string.h   basic_string.tcc   locale_classes.h   stringfwd.h   basic_ios.tcc   exception   functexcept.h   debug.h   predefined_ops.h   new_allocator.h   locale.h   atomic_word.h   atomicity.h   <built-in>    new     ���  ��� ���~X  М� J�J�~<�f�~�   �� �  @�� ��<�}= �%  Н�   ��    �� JO�   �� JO�  @��X����~�u�~Xz<Pz<�J�~X��  ���t	< 4� L�X��.� <�Xzf� t�.� <v��C.=<�<Og?X��.� <�XO� f�CX:X�  p���l�.� ���vJ
<v<
�x��.� <�<Og� X��.� <�<O� f��X� X�  `���B�l��zfBX�~.�<�Xzf� ��.� <�<Og� X��.� <�XO� f��X� X�  `�����@<2<Nf2<X�~.�<�~Xzf���~.�<�~<Og�X��~.�<�~XO�f��~X�X�  P���  ����� <�= �$  �-X�+i K��?� �z<��� X  ���XM �� �~J ���d�}<�<�}Xzf��  �� j8<juqtXq�f
.v<Xz<����~J���}�����}<�<�}Xzfx�s�XtX�.b<<OgdX�.f<XOef�Xdt  P��	fw<<	fu���Z� J�J��~J���~��<�}<�<�}Xzf��J	�~.�.	�~<�<�}��i.<oXzf��z.Bu<Og[
XyJZ�v.
<qXO	fx�|  ���
fv<<
fu� ��.�~fK�~.�<�~Xzf����~J���~��X�}<�<�}Xzf6�w�\.$<W<Og&X�X.(<SXO'f�U`WJ&t  ��   ��XK�.�|t�J�}��jJX�ȑ�y%  ���=  ��� 
 Ш�<L�tf
�~��<�|<�J�|fnXJ
�~<�t��y� 
 P�� La�
!t 
 p�� L_
yJ5t.
C 
 ��� � X � � �t j
 � X 
 ���J
�|J�.
�|t 
  ���J
�|J�.
�|t   �� lz<<Bu��;gt.�Ʉ���~t��~J���}��<�|J=I/� <Bzf�&�| Y� .�<� XzfI� fK�f�}.	����� f�|J�J_�}�Z��<�}�	���f� J�|J�J_�}�Z� .�<� Xzf���}<�<�}XzfY��%�|<�.�|<�f��|tKI� ��|f�Jg�|J�� �;=Ց-=�y.���z*�9.G<4<OgIX�5.K<0XOJf�U`4tIt   ��<�  @��v��  `����  ���X�	�}J���}�}.�<�}Xzf��  ��Xp�	�}J���p��}.�<�}Xzf��  @��Xu�	�}J��	�u��}.�<�}Xzf��  ��>i9<?u�h����X�J�n�f� .�<� Xzf����~J���}��J�|<�.�|<�f��|�Y� ��}<�<�}Xzf���J�;=�y1J�� .�<� <Og�X
XytZ�� .�<� XO�f� ��t  ���  ��� �lXt�   ��   �>i9<?u�h����X�J�n�f� .�<� Xzf����~J���}��J�|<�.�|<�f��|�Y� ��}<�<�}Xzf���J�;=�y1J�� .�<� <Og�X
XytZ�� .�<� XO�f� ��t   ��  0��  @��  P�>����h����X�o��X�n�f� .�<� Xzf����~J���}����|<�.�|<�f��|�Y� ��}<�<�}Xzf���J�;=�y1J�� .�<� <Og�X
XytZ�� .�<� XO�f� ��t  p��  ��>��G?g�h����X�J�n�f� .�<� Xzf����~J���}����|<�.�|<�f��|�Y� ��}<�<�}Xzf���J�;=�y1J�� .�<� <Og�X
XytZ�� .�<� XO�f� ��t  ���  ��>��G?g�h����X�J�n�f� .�<� Xzf����~J���}����|<�.�|<�f��|�Y� ��}<�<�}Xzf���J�;=�y1J�� .�<� <Og�X
XytZ�� .�<� XO�f� ��t  к�  �>i9<i+?Y�h����X�J�m�f� .�<� Xzf����~J���}����|<�.�|<�f��|�Y� ��}<�<�}Xzf���J�;=�y1J�� .�<� <Og�X
XytZ�� .�<� XO�f� ��t  ��   ��@�   �>i9<?u�h����X�J�m"f� .�<� Xzf����~J���}����|<�.�|<�f��|�Y� ��}<�<�}Xzf���J�;=�y1J�� .�<� <Og�X
XytZ�� .�<� XO�f� ��t  0��  @�>i9<?u�h����X�J�m�f� .�<� Xzf����~J���}��J�|<�.�|<�f��|�Y� ��}<�<�}Xzf���J�;=�y1J�� .�<� <Og�X
XytZ�� .�<� XO�f� ��t  P�� V   Q  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include/sys /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  locale_facets.h   stdio_sync_filebuf.h   streambuf   postypes.h   char_traits.h   basic_string.h   basic_ios.h   c++config.h   allocator.h   cwchar   clocale   basic_string.tcc   ios_base.h   cstdio   c++io.h   ostream_insert.h   debug.h   predefined_ops.h   new_allocator.h   cpp_type_traits.h   stddef.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   types.h   file.h 	  wchar.h 	  locale.h 	  functexcept.h   atomic_word.h   stdio.h 	  new 
  <built-in>      ���  `�7�J  ��7J�J�~�  ��� J� J��>  ��� J� J���  ��� J�� X��vu�[  0��  @��4zX<�].#�3�=[
  ���<  ���X��� t��Hv   ��<�=XM�3<E �x<`  p��XO�4JLX*�S<-�
 w�	X&   ���l<�f�   ��XL�m.�|t�J���p��y%  ��� J�J�|9=   ��     5  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  istream.cc   char_traits.h   streambuf   basic_ios.h   ios_base.h   ctype_inline.h   basic_string.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   c++config.h   cwchar   clocale   allocator.h   basic_string.tcc   locale_classes.h   stringfwd.h   ctype_base.h   istream   istream.tcc   basic_ios.tcc   postypes.h   stl_algobase.h   locale_classes.tcc   debug.h   predefined_ops.h   new_allocator.h   exception 	  locale.h   atomic_word.h   <built-in>    ctype.h     �&i9<gv����~���L�j<�~�:h;=-=�Y:����~��.�~<�t�~.�.���zXZ�<�<�|<�<�z<�<Lf�~��� .�<=XO��I�<�ug� t@<..R<4Xz<T�Me�Z� <�X0�����|<�.�}t� .�~<�<�~�=�J�J�~fLJ�~f�<m�h��~���m2�}�2Ȓ� .�<� <Og�Xt�� ��t   �� ��=;u�{�f�~J�L�jf!<_J�~�eg���� ���� .� <�~<�J�z<�<�z.�.�z<�<�~.�<Lf�~<eg"Jgh�j�)<^��=Ite��f�~.�<�f�~�Lt7��~�� p�ev���X�~�h���Zf&<`Xzf��m<�~�kf<fXOgX�gf<bXOf��kXt   ��
fv<
<���f�|<V��X�|��<�|X1� f�<� L�Vfj. �~J �< �~.��䱏>:���<� <�<��0:� J%.���{<� <�<�<�|X�<�|<�f� f@<f�<�J�|<=�X�|����f� <�XO� �[�fBz<� �p��<�|<=�X�|��f��� <�t�uM#t�-<S<� �� �=I�  ���~fL�V<�~�.qּuM�!fY.! l-t;��!X*1b�fq�f\�$fb���_���m<h�JX5<,���� ��~"7��f� <�XOg� t�RtJX� t   ��fu<<�9���~fBz<�<���<�z.�.�w��f�<�w V��X�|X�<�|X � � (f X< (L� �< �|� �< �~.���e"��~<�<�~<��&:�J;/���|<>�<�|X�<�|<]fof<fZ�<�}<�.�}f�<�}<�.�}��~���� <�t�uM#t�-<S<� ����X�<=��yf2X�X� �y����~f�Z��<�J�}<�.�}��}�.qּuM�!fY.! l-t;��!X*1b�fq�f\�$fb���_���h�]��
t<� �Y�(��~f�<�~XOg�Xu<8�w��Z��~f�<�~XO�f`�~��t  ���ft<<<����X�}f�<�}Xz<�����<�z.�.�w�� ��<�x<Z�L�j<!._.� �=sv��� �X�<����|<>�.�|.�<�|<Lf� <Z��~"
.�X�<=;=��y�2X�X��<�J�~f1(�<��h����v<
t<���f�X�f��m���xt��}f�<�}XOg���Z��}f�<�}XO�f�}f�t y|   �  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  locale_facets.h   locale_facets_nonio.h   locale_facets_nonio.tcc   messages_members.h   locale_classes.tcc   locale_classes.h   time_members.h   codecvt.h   basic_string.h   atomicity.h   char_traits.h   c++locale.h   ctype_inline.h   ios_base.h   streambuf_iterator.h   streambuf   locale_facets.tcc   locale-inst.cc   locale.h   clocale   cwchar   cpp_type_traits.h   stl_iterator_base_types.h   stddef.h   c++config.h   allocator.h   basic_string.tcc   stringfwd.h   ctype_base.h   ctime   postypes.h   stl_algobase.h   stl_iterator_base_funcs.h   functexcept.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   type_traits.h   debug.h 	  predefined_ops.h   new_allocator.h   stl_iterator.h   atomic_word.h   time.h   new 
  ctype.h   <built-in>      ���  ���  ���	  ���	  ���	  ���	IK  ���	IK  ��	   ��	  0��	  @��	IK  `��	IK  ���
  ���
  ���  ���  ���  ���  ��?  ���    �� N*N Y e = -P  0��  @��  P��  `��  p��P  ���K  ���VJ  ���  ����~J  ���	KIK  ���	KIK   ��	KIK  P��	KIK  ���	KIK  ���	KIK  ���	KIK  ��	KIK  @��KIK  p��KIK  ���KIK  ���JLQyf0 t� t� t� t�  @��JLQyf0 t� t� t� t�  ���JLPzf0 t� t� t�  ��J	J  0��J	J  P��
J  ���
J  ���J  ���J  ��JR  0��J  `��J  ���J  ���JP  ���JK  ��JVJ*�  @��J  p��J�~J��  ���J��  ��:X= %  �:JK  0��K  @��JK  p��X= %  ��� X>@bY �� t��;=   �� JP  @��  P��J 	 ���
�~J=	�<
�~.	�<5��  ���	�f�s<<	�<�s'>	�<�s�0��� t��� .��/�	� tCf=tCfStx�O=p<	� �Cf=�CfS�y<	� �Cf  ����g�;/ǟ  0��X�<� t�f  p��X=>  ���X�<� ��.  ��	�f�s<<	� ��f�t�>,Z:>>
t˅;==Y�;/��c�/	:XI.	�<�<=;=��y<	2J�.�v<
t<O	5�C<=<C<tw&	;XCf=�CXv���  ��:1U!�r0	�O9.i���;/��OyX5Y�  ���t��L�����s   �2uI�u8�o�ztg��M,Sf2�N<2.T.�!Y� 	Y�!<e�q�n��\�$�1b�k�t�  P���{ �.�{J�<�{<�.�{��<�{<�<W  ����{ �.�{J�<�{<�.�{f�<�{<�<gW  ����{ �.�{J�<�{<�.�{��<�{<�<s  @��K���~t
  p��K���~t
  ���J����~f#   ��J����~f#  `��J����~f#  ���J����~f#   ��K���~f  P��<�� ���(  ���<�� ���(  ����{ �.�{J�<�{<�.�{��<�{<�<W  @���{ �.�{J�<�{<�.�{f�<�{<�<gW  ����{ �.�{J�<�{<�.�{��<�{<�<s  ���K���~t
  ��K���~t
  @��J����~f#  ���J����~f#   ��J����~f#  `��J����~f#  ���K���~f  ���<�� ���(  @��<�� ���(  ����{�J�{J�J�{��<�{��<^   ���{�J�{J�J�{��<�{��<^  ���
�x �.�x��<�x<�.�{��f��:h�}��< K �RF=��v��}  ���
�x �.�x��<�x<�.�{��f��:h�}��< K �RF=��v��}  P��
�x�J�xJ�J�xf�f  p��J�2  ���J�2  ����v�	J�vJ�	J�vf�	f  ��J�4  P��J�,  ����u �
.�uJ�
<�u<�
.�u��
<�u<�
<;  ����u �
.�uJ�
<�u<�
.�uf�
<�u<�
<g;  0���u �
.�uJ�
<�u<�
.�u��
<�u<�
<I  ���K� ��t
  ���K� ��t
  ���J�� ��f#  @��J�� ��f#  ���J�� ��f#   ���v�	J�vJ�	J�v��	<�v��	<)  `���t �.�t��<�t<�
.�u��
f��:h�~��< K �Rb/��v��~  0���s�J�sJ�J�sf�f  P��J�,  ���J�,  ���J�,  ��J�,  P��J�,  ����q�J�qJ�J�qf�f  ���KW�#  ���J�*  0��J�.  p��J�&  ��)� �}.�J�}<�<�}.���}fY;=��  �1� �}.�J�}<�<�}.�f�}fhY;=��  p�9� �}.���}<�f�}.���}f|?�pȻ��rX�g ��	  P����
  p����
  �����
  ���  �����
  ����������
  0 ��������
  � �������������  �������������  �� ��~J�J�~J���~<���~<�  P��}�J�}J�J�}f�f  p�LV�-  ���|�J�|J�J�|f�f  ��lJlJJkff  ��K   �J�,  @�J�,  ��J�,  ��J�,   �J�,  @��}�J�}J�J�}f�f  `)�.�}.�<�}J�J�}.�f�}f�  �.�.�}.�<�}J�J�}.�f�}f�  ��K  �4L   �J�   0�K  @�g  P�	�sJ�f  `� iU<=�:h = �P��x�  ��iU<=�:h = �P��x�  ���~.�.�~<�J�~J�.�~f�f� �  ���~ �.�~<�J�~J�.�~f�f�  ��L   �J�  0�K  @��| �.�|��<�|<�.�~f�f�X�~<�<Vh � �P���x��~  ��>�K;/;= .w�zJ Z  @	���|���g<m��~J���~.�����~J���~.�����~J���~.��.l[���~X���z��.�xJ���� .�X�K��K��.�~�||�~�>   �	JwX�~��t� � �z $�� ��.��J�Y�� i��z�����<v�Y ���z��.�z.�X���}f�X�{�L��t��L�4fL��<��{f�$�{��~��� ��~��<�~\�J�~��f�~.��t�z.�   �t�|��<jH�3��x��V� J�.���xJ�t��x��.LX4��~����~�#� �3X�~�  ��>�K;/;= .w�zJ Z  ��>�K;/;= .w�zJ Z   �>�K;/;= .w�zJ Z  p� �>L��� .	�t�D�<�|<=f�~<	�<�~f�;=�<� � �r�	 �� �~<	 �< C<�~�=;= f  �<� �	�s��<�|<C<�~X	�<�~f�;=�<� � �r�	 �� �~<	 �< C<�~��f� �	�s��<�|<C<�~X	�<�~f�;=�<� � �r�	 �� �~<	 �< C<�~��f� ��rt�<� ��rt>���yJ=��O��.�~5�y<�����.�x+���;=�y��<��;=�y��<�y� ��G�s�,� � � �
�r`=	�<
�~.	�<j
�~�=	�<
�~.	�<j�~"�	 �X Cf��_�s $t �Y t�_B!t	 � Cf =� Cf  ��>�K;/;= .w�zJ Z  �>�K;/;= .w�zJ Z  `�>�K;/;= .w�zJ Z  �� �>M���.�wt�<���wt�<���vf�<��	�x��<�|<C<�~X	�<�~f�;=�<�� �w�	 �� �~<	 �< C<�~�=;= f  �<��	�x��<�|<C<�~X	�<�~f�;=�<�� �w�	 �� �~<	 �< C<�~��f��	�x��<�|<C<�~X	�<�~f�;=�<�� �w�	 �� �~<	 �< C<�~��f��	�x��<�|<C<�~X	�<�~f�;=�<�� �w�	 �� �~<	 �< C<�~��f� � �wf �<� ��vf>���yJ=��OL���x���;=�y��<�y� �J� L�� o�� o� � s��?���s��x�ss$t � �Y t� t�	 �X Cf�~s!"�	 �X Cf��^�ss$J	 �* Cf =# Cf<  @ �>�K;/;= .w�zJ Z  � � �>M���.�wt�<���wt�<���vf�<��	�x��<�|<C<�~X	�<�~f�;=�<�� �w�	 �� �~<	 �< C<�~�=;= f  �<��	�x��<�|<C<�~X	�<�~f�;=�<�� �w�	 �� �~<	 �< C<�~��f��	�x��<�|<C<�~X	�<�~f�;=�<�� �w�	 �� �~<	 �< C<�~��f��	�x��<�|<C<�~X	�<�~f�;=�<�� �w�	 �� �~<	 �< C<�~��f� � �wf �<� ��vf>���yJ=��OL���x���;=�y��<�y� �J� L�� o�� o� � s��?���s��x�ss$t � �Y t� t�	 �X Cf�~s!"�	 �X Cf��^�ss$J	 �* Cf =# Cf<   (�>�K;/;= .w�zJ Z  p(�>�K;/;= .w�zJ Z  �(�>�K;/;= .w�zJ Z  )�	��|t�f��}��t�}.g�J-g�0rg��xt�.�xt4n<.���~�q?�~��r.us�} �6  �*�>�K;/;= .w�zJ Z   +�>�K;/;= .w�zJ Z  P+�>�K;/;= .w�zJ Z  �+� L�M91U? . t �  �+� L�M91U? . t �  @,� L�M91U? . t �  �,� L�M91U? . t �  �,� L�M91U? . t �  0-� L�M91U? . t �  �-� L�M91U? . t �  �-� L�M91U? . t �   .� L�M91U? . t �  p.� L�M91U? . t �  �.� L�M91U? . t �  /� L�M91U? . t �  `/� L�M91U? . t �  �/�	3)��|�2/ � 7.�xJR/�/;�d�YIY " �G'� & ��� k �yJ  `1�t| M c 1 + 1 � �z. �< i / �z. �� v / vJ w ^ /   2�X��K  @2�����}f� �}<�}X�t�}<u=;=	�.�X�Y;g�}<�<�}<��%:K�.�	�~f�t�T@Y-=h0:h�	�.�z<	�.�|<�<�z�	�.�z<	�~J�<	�~<u� 	�~X�<	�~<u� 	�.�}<nJ���x�j	�J�|<	�<�|<�%�|<�<�|f�<�|<���|<�< � 2	 �~� �t v : h > , Z !� _J !<d�t r�%�g	�~��<�~<�	���y�	�X�w�f�~<	�C<=�Cf�X�<� <�t!��=;=	�<�}<>=-=�}.�<A�}<���� <�Je��uM!6�S�� ��(�.y�	�f�|��	�X �|�k���;=�| $.1n�tY�^!�; ;���wt	�bt�\t$�qt�Lf���t�yu�y<C�f	���z"	(JiCf=�Cf�~t�U��  `:�����}f� �}<�}X�t�}<u=;=	�.�X�Y;g�}<�<�}<��%:K�.�	�~f�t�T@Y-=h0:h�	�.�z<	�.�|<�<�z�	�.�z<	�~J�<	�~<u� 	�~X�<	�~<u� 	�.�}<nJ���x�j	�J�|<	�<�|<�%�|<�<�|f�<�|<���|<�< � 2	 �~� �t v : h > , Z !� _J !<d�t r�%�g	�~��<�~<�	���y�	�X�w�f�~<	�C<=�Cf�X�<� <�t!��=;=	�<�}<>=-=�}.�<A�}<���� <�Je��uM!6�S�� ��(�.y�	�f�|��	�X �|�k���;=�| $.1n�tY�^!�; ;���wt	�bt�\t$�qt�Lf���t�yu�y<C�f	���z"	(JiCf=�Cf�~t�U��  �B�� f�<<� ���� X � : h	 �}� �<	 �}< <u� �����|< e K	 �}� �<	 �}< C<��� I��-=�}��f�}<�.
�y�=	�<
�~.	�<j4�Cf��  `D�NT� . 5 ; =!  �D�	t�F�w��<�w.�X�/�x����x.�X�xJ�J�xJ���xt� �|<�<�}f�t�}.�f��}X�JpJ�/Y�xf�X�x.j��xt��M;V=�}����}����}����} ���}�%   G�X��W�/  PG�NT� O r 0 Y - ,.K�zX�t�zX�J�z.�X # / ; d 0 d u� / ; d 0 r   H���y<�X�y�u=;=�.Bztl�y<�.�y<�<�y<�<�=;�N91F\9?����M�;K�=!�}.�}����~�?�~���^ r��;K->;KI���>�=;@;9=[9>t��y����z<� �	t�yf�<�t:{y<C�<�yt��?U  K���xX�<�x.�<1s/;=(�K;=�w�!=�X � > : k�[�y��J�yJ�J�y<�~��<�|<�t�wf�X�y����~����~�9?�fPz<B af > : k�y��J�}t�f�~�9?G���~���~�?�~f���z<;� �	t�t@����~Ȓ�?U   N�JK)  @N�X�� �~�4  �N���y<�X�y�u=;=��Bzt�
<�yf�X�y<�<�828@�?8Y[��M�;KW=u�}.�}��f�~�?�~���P��;�->;KIPF�fh��;@;:[9>�y����	t�y@�zf{y<C�<�yt��?U  `Q�JL)  �Q�	t�w�x���W�{f�<��  R�X�� �~�4  �R�xT@ � � � 1 q 1 G.K;/�zX�t�zX�J�zJ�X � = � , u� g � 1 G 1 G  �S���yf�X�ytu=;=��Bztl�y��<�y<�<� � � � 9 1 F Y ?f��.M�;K�=!�}X�}��J�~�?�~���^Jr�;K->;KI&p2f���;@;:[9>tt�y����z<� �	t�yf�<�t:{y<C�<�yt��?U  �V�JL-   W�t=� �~X,  �W���yf�X�ytu=;=�.z<BzJl
<�yf�<�y<�<�8282=?8Y[��M�;KW=u�}.�}��f�~�?�~���P��;�->;KI"�����;@;:[9>�y����z<� �	t�yf�<�t:{y<C�<�yt��?U  PZ�JL-  �Z�t>� �~X,   [*�>�/�tf���t�yu-=��w��U��  0\*�>�/�tf���t�yu-=��w��U��  `]4�>�/�uf���	t�t@-= X C �x��U��  `^�
fvX<�} �<CyJ��	<w<	.w<	<taffɄVL�>�zfBi�~�̈́��yJ� �;Yl�M�;Ks=Y�|f�}t�f�~.9?�~���Y� � X �ut.1;6>:"�>H��~�!��~.��=�Y�~�  @a�JL/  �a�
fvX<�}��<yJ��	<w<	.w<	<taffɄVL�>�zfBi�~�̈́��yJ� �;Yl�M�;Ks=Y�|f�}t�f�~.9?�~���Y � X �ut.1;6>:"�>H��~�!��~.��=�Y�~�  `d�	JM3  �d�JN�	X��LX�<A� �~��itX  e�X	����v�� LX�<�tLX�<rX���~���.�~��p��   f��~��f��z �<�zJ�t�z<�f�z��f�-=�y����. �" � � �������z.�f�zX���z.�< L �z< �X�y������}f�tu�z����Yb2*0=;/�z��X�z<���L��<�z<�<1z<wJ��y�v����zX�<=e�z<���z.�.�z���w��{�~��x�� � �yJ �t �y< �X�y�v���;  i��zf�<�~<�f��zX�<�zX���0s �yX��� t�.���y����% pL�;�v�;==w<6YwX.�y������}f�t�z.LX�<Bz<� L��<�X� ��yX�f�-=�z.L��<���~��xt� t � �< ���zf�~����~��G��<�y.� �y.�X�. �~' �� ������yX�<�yfL��� * �z< �� �z< �< ;�  ��y.��s�s  m��}t�t�}��<��y��=;KK���n�������<�y�u��l��xքV� J�.���xJ��Y�x��.LX4��~����~�#� �3X�~�  0o��}��t�}��<��y��geKK��������dȟ�����������<�y���l��xքV� J�.���xJ��Y�xX�.LX4��~����~�#� �3X�~�   r�� t��g;3*�}X���}.�� �|<��� ��.������}.����}��.�}�;��2�}��~��x��� ��X��L��<�����z����-=�z��J�z<����z��X�}�L��<�!K�}����}��.�!��{�L��J�|����}f�J!�yJ���~���� �:�}��|��<��@�{����~X�{XfJ���~X�{X����Z��{'����{�����y�!�=J�|@�<�|�ɟ���������o��JYp��|:�uu���tf�JY�{�����{^�t � ��z��<�AJ�zf�<�AJ�V�{]�<q�Kr�v�Ks�!�t<!�7!�z<K� �]��|4�uu��������]��uu���� ��~��&�~t!��f��V�{<��K�{f�J�zf  @�t�}��<�yf�<�y/�X�yJhV� J�.���yJ�t��z�LX4��~����~��� f3��~�  `��t�}��<�yf�<�y/�X�yJhV� J�.���xJ�t��z�LX4��~����~��� f3��~�  ������{f�	�x<Dw<	<xJD J �	 � < �tg	� f�t�=q?W=;=\� ) �~� � ���� ��.� � ���]�'.�� t�.2�L��� �c�	5��<�<=��yX	2X�<��<�����}f\.$t�� f�X�L��<.XL�	�J�|<��0f�Ȅ	U�+<	U<C<=�Cf� ��~���U< � J � � xJ ��� .�GM��	�J�|<h0K	�X�|< f$	jf<�h�<:	Yu���v<�	<�v<�t�|<w	���z<	�< �z�	 �< �z< � f(%L��<Bz<���L��<�~f���~�'��� f�X��L��<�.L��<Bz<�.L��<8��I� � ��	���zJ�~.��KM�t�-<S<�!�h"�_�����~�����~��	�
t<� Xz#���}f���~�����~�����~�� SJ=- p���� t�.��.� ��<� <� �D��.�~�\xtv� f�X��L��<X��JLX�<SJ���X�}f 6t� <��~�����~��G���~���� �+����� Jz�1� �� ��~W� ��~�� ��<� <������ � 
��  � � �� � � �< � <��~X���~f�<�~X���X�}f �tf�~�� ��<� <������ � � ��~���X	T�Cf=�Cf  0�����{f�	�x<Dw<	<xJD J �	 � < �tg	� f�t�=q?W=;=\� ) �~� � ���� ��.� � ���]�'.�� t�.2�L��� �c�	5��<�<=��yX	2X�<��<�����}f\.$t�� f�X�L��<.XL�	�J�|<��0f�Ȅ	U�+<	U<C<=�Cf� ��~���U< � J � � xJ ��� .�GM��	�J�|<h0K	�X�|< f$	jf<�h�<:	Yu���v<�	<�v<�t�|<w	���z<	�< �z�	 �< �z< � f(%L��<Bz<���L��<�~f���~�'��� f�X��L��<�.L��<Bz<�.L��<8��I� � ��	���zJ�~.��KM�t�-<S<�!�h"�_�����~�����~��	�
t<� Xz#���}f���~�����~�����~�� SJ=- p���� t�.��.� ��<� <� �D��.�~�\xtv� f�X��L��<X��JLX�<SJ���X�}f 6t� <��~�����~��G���~���� �+����� Jz�1� �� ��~W� ��~�� ��<� <������ � 
��  � � �� � � �< � <��~X���~f�<�~X���X�}f �tf�~�� ��<� <������ � � ��~���X	T�Cf=�Cf  ���k7AE	��� t . %XK	�~<�<	�XDC<�� T
�}�=	�<
�~.	�<24Cf  Н����}<�<�}<iU	�.� t X	 �. � <	 �< �}<O	�f� <	�~<�f	�~X�f w�	�0�|��<�|<JuhJ�f�L���~�
�y�=	�<
�~.	�<j���| �X	�{ Cf  ���
fv.�<�{f6�R�.XR<� 	� .�tj�� 	�v��z �X�����}<�t�~fL��<Bz<� ��.� �	(�:<w3�	B�><	�<� ��~<� X X	���y�	�<�y<�����}<�t�~fL��<Bz<� J�.4���� �,<T. f y< Qg	 �X �y�	 �< �z< �J'Ȯ� f�X��L��<� X����U�� .L��< " s	���z�� ��~�$t����~�����~��xt� �^�M�7  J�n�%<�	�<�z<	�<�z�	�J�z<�~X�����}<�t�~fL��<Bz<� J�.���~����~f�<�	���y�	�<�zt�~t'��� f�J��L��<�X��	���|<	�t�z$  X ��	���y�	�<�y<�t���}f� t� .�~���W<*. Xy� ` IK ��	�X�{<	�f � �z<��~�$t����~�����~�$t���~�����~����x.	U.�����a<.= ��X J X��T�1<OJ�����}<�t�~fL��<Bz<� ��.
�	� ':< �~� IK ��	�X�y<	�f�y���� �U�[�	�t:<	���{#L��<^C�	�$�y�	�<�y<OJ'�� � J�~�\<$t�t1�~�����~���<���~����	��� <�.� .�{%Cf  ���k7	�|<���0�|��d� J�.���{f�f	�|��<	�|<C<���}LX�<�X�~����~�\xt� J
�~ =	�<
�~.	�<2� .�~�	� Cf  ��k7	�|<���0�{��d� J�.���{f�f	�|��<	�|<C<���}LX�<�X�~����~�\xt� J
�~ =	�<
�~.	�<2� .�~�	� Cf  `��k7	�|<���0�{��d� J�.���{f�f	�|��<	�|<C<���|LX�<�X�~����~�\xt� J
�~ =	�<
�~.	�<2� .�~�	� Cf  Ю���<�}<�}��<x<D�}t�< X �~. �� �~X �<�}f���f� <= � s ��~�v�� ���+�_Js/� � j	 �~. �tmg-�ihH>��֜�&�sf�}��<�}X�����}<�t�~fL��<Bz<� ��.��c�	�~f�<t���|f�f	�}f�<	�}<�X	�}X�f	���|	�<�|<M�	�}��< �����]���u�sf�K�/H�}.'��� f�X��L��<�X�}����L��<�J�q��~�$t����~�����~��G����< ���~��.�0�\K�I-�|.�����}<�t�~fL��<Bz<� ��.���|t�<�|X'J�� f�J�XL��<��	���|.�~ �~�$t�t1�~�� ������~��~�����~�����}���� �� J ��
� � ���s�}������}f� t�� e)�M�}����~t�f�f�3�~�.�� X�XoN	��Cf  ���JL/  ��J����~&9  `��tN��7IK��|J�<=�|����|���� <�<V�g:YY���|ȼ�� ��X���|����K��K���|��J�|<�t���}f�� � g � cf�!. f�Wui ��}fL��<�f�Xn ��}fLX�<zJ�<LX�<���~�$x�� �3��~�\��� ��-=y<L,>�|.�����u�}��~�\� x �  м���<�}<�}��<x<D�}t�< X �~. �� �~X �<�}f���f� <= � s ��~�v�� ���+�_Js/� � j	 �~. �tn�hH>��֜�&�sf�}��<�}X�����}<�t�~fL��<Bz<� ��.��c�	�~f�<t���|f�f	�}f�<	�}<�X	�}X�f	�t�|	�<�|<M�	�}��<A*]���u�sf�Y�/H�}.'��� f�X��L��<�X�}����L��<���q��~�$t����~�����~��G����< ���~��.�0�jY�I-�|.�����}<�t�~fL��<Bz<� ��.���|�<�|X'J�� f�J�XL��<��	���|.�~ �~�$t�t1�~�� ���I��~����l��~?�~�����}���� �� J ��
� � ���s�}������}f� t�� e)�M�}����~t�f�f�3�~�.�� X�XoN	��Cf  ���JL/  ���J����~&9  p����<�}<�}��<x<D�}t�< X �~. �� �~X �<�}f���f� <= � s ��~�v�� ���+�_Js/� � j	 �~. �tn�hH>��֜�&�sf�}��<�}X�����}<�t�~fL��<Bz<� ��.��c�	�~f�<t���|f�f	�}f�<	�}<�X	�}X�f	�t�|	�<�|<M�	�}��<A*]���u�sf�K�/H�}.'��� f�X��L��<�X�}����LX�<���q��~�$t����~�����~��G����< ���~��.�0�\K�I-�|.�����}<�t�~fL��<Bz<� ��.���|��<�|X'J�� f�J�XL��<��	���|.�~ �~�$t�t1�~�� ���I��~����l��~1�~�����}���� �� J ��
� � ���s�}������}f� t�� e)�M�}����~t�f�f�3�~�.�� X�XoN	��Cf  0��JL/  p��J����~&9  �����<�}<�}��<x<D�}t�< X �~. �� �~X �<�}f���f� <= � s ��~�v�� ���+�_Js/� � j	 �~. �tn�hH>��֜�&�sf�}��<�}X�����}<�t�~fL��<Bz<� ��.��c�	�~f�<t���|f�f	�}f�<	�}<�X	�}X�f	�t�|	�<�|<M�	�}��<A*]���u�sf�K�/H�}.'��� f�X��L��<�X�}����LX�<���q��~�$t����~�����~��G����< ���~��.�0�\K�I-�|.�����}<�t�~fL��<Bz<� ��.���|��<�|X'J�� f�J�XL��<��	���|.�~ �~�$t�t1�~�� ���I��~����l��~1�~�����}���� �� J ��
� � ���s�}������}f� t�� e)�M�}����~t�f�f�3�~�.�� X�XoN	��Cf  ���JL/  ���f��z�\�f$�~��</�-=	  `��J����~&9  �����<�}<�}��<�}��<�}<�< . �~. �� �~X �<�}f���f� . � I ��~�v�� ���+�_Js/J � j	 �~. �tm " � 9 i >�+ f��~��X�1;�;=@u;�4gI�|f�����}<�t�~fL��<Bz<� ��.����	�~f�<t���|f�f	�}f�<	�}<�X	�}X�fP	���|	�<�|<�M�	�}��<��s��}��<�|X'��� f�J��L��<�X�|�����	���|.�~ �~�$t����~������&�s��}��<�}X�����}<�t�~fL��<Bz<� J�.���}��\�.�����q L��<�u;�%gI�}<�<�}<'��� f�X��L��<��q��~�$t�t1�~�����~�� ���I��~����hL:j��~`�~�����}���� �� J ��
� � X�s�}������}f� t�� e��MF�}f���~t�.� ��~����~�.�� ��.oN	��Cf  ���JL/   ��J����~&9  ���fnX<�<�}<�}��<�}<�<�}<�< . �~� �� �~X �<�}f���f� <= � s ��~�v�� ���+�_Js/� � @	 �~. �tni9i>H>�����&�sf�}��<�}J�����}<�t�~fL��<Bz<� ��.��c�	�~f�<t=;�f�|f�f	�}f�<	�}<�X	�}X�f	���|	�<�|<�M�	�}��<A�]���=e�u�s��-Y;u-=�/$�}.�</I�}f'��� f�X��L��<�X�}����LX�<���~��~�$t����~�����~����YKI�|f�����}<�t�~fL��<Bz<� J�.���|����< ���~��.�190���-Y;u-=�/�|1�<�|J'��� f�J��L��<�f	���|.�~ �~�$t����~�� ���I��~����l��~Z�~�����}���� �< J ��
X � ���s�}������}f� t�� ef�M8�}����~t�<�����~�.�� ��XoN	��Cf  P��JL/  ���J����~&9  ���������������n������	��w� N   �  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  allocator.h   c++config.h   debug.h   predefined_ops.h   new_allocator.h   cpp_type_traits.h   <built-in>    new     ��    ��   0��   @��   P��   `��     z  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  locale_facets.h   ctype.cc   locale.h   clocale   cwchar   char_traits.h   stddef.h   c++config.h   allocator.h   basic_string.h   basic_string.tcc   locale_classes.h   stringfwd.h   ctype_base.h   ctime   stl_iterator_base_types.h   cstdlib   cstring   ctype_inline.h   c++locale.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   debug.h   predefined_ops.h   new_allocator.h 	  stl_iterator.h   cpp_type_traits.h   atomic_word.h   time.h   stdlib.h   string.h   new 
  <built-in>      ���  ���  p�4X>dh�� J�Aa  ��4JO  ���J��  ���J��   �� 0,� ? ;��f�w0;u	.v����wXMr�
�   �� 0,� ? ;����x*:L/Kz�    g  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include/sys /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  ios_init.cc   streambuf   stdio_sync_filebuf.h   basic_ios.h   ostream   istream   ios_base.h   atomicity.h   stddef.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   types.h   file.h   wchar.h   char_traits.h   c++config.h 	  cwchar   clocale   ostream.tcc   cstdio   c++io.h 	  basic_ios.tcc   fstream   iosfwd   debug.h 
  predefined_ops.h   new_allocator.h   exception   locale.h   atomic_word.h 	  stdio.h   new   <built-in>      ��� {d�t�|P	f�f�|t�<�|K
f�f�|t�<vK�}t���}X���}@���}����}@��X�}����}@���}����}@���~����~�/t�X�  ��� uY<t.f  ��� HY;<E<;f.h�f���+�  P��wqC��g<t.f� f]<#Xo@����s� }   %  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/tr1 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/MXlibraries/include/sys  stdio_filebuf.h   fstream   streambuf   ropeimpl.h   stl_iterator_base_types.h   cstdlib   new   c++config.h   allocator.h   cwchar   <built-in>    tuple   functional   cstdio   char_traits.h   postypes.h   clocale   ios_base.h   functexcept.h   basic_file.h   c++io.h   fstream.tcc   cpp_type_traits.h   debug.h   predefined_ops.h   new_allocator.h   memory   rope   algorithm   functional   ext-inst.cc   stddef.h 	  stdint.h 
  kernel.h 
  fs.h 
  ipc.h 
  kernquery.h 
  stdlib.h   types.h   file.h   wchar.h   gthr-default.h   stdio.h   locale.h     ��� X� <j��j<�<� f�j�  �� JK  0��
J�>JJd�=0x���s�vX/  ��� J  ��� �g":Z:h� ���	JzX=:==�f�}<I>�J�Qt==�}<t�  p���h":Z:h� ���	JzX=:==�f�~<I>�J�Qt==�}<t�   �� 
  0�� 
 �   �  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext  streambuf.cc   streambuf   char_traits.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   cwchar   clocale   c++config.h   postypes.h   locale.h   debug.h   predefined_ops.h   new_allocator.h   atomicity.h   <built-in>      @�&tMGM�fL��~<�Y�X�|��<�z</�J�}���.Z� .�|��<�J�~fLJ���~f�<�}X�|�.h�+f�}X�.�}J �   /  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  sstream   streambuf   sstream.tcc   char_traits.h   basic_string.h   atomicity.h   basic_ios.h   ios_base.h   stl_algobase.h   postypes.h   istream   ostream   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   cpp_type_traits.h   stl_iterator_base_types.h   c++config.h   cwchar   clocale   allocator.h   basic_string.tcc   basic_ios.tcc   stl_iterator_base_funcs.h   debug.h   predefined_ops.h   new_allocator.h   stl_iterator.h   type_traits.h   exception   locale.h   atomic_word.h   new   <built-in>      `��M� ����}X*  ���O� ����J��}�  ��,<�]�X$<�~.���|<�.�|</X���~<�.�|<e�  ����~J=�<�~.�<2�  P�?X�J�~<�fC<V��~ =�<�~.�<2  ��?X�J�~<�fC<V��~ =�<�~.�<2  ��X�~J�<�|��tC<V�� ��<� f���|=�<�~.�<2�.  ���XTJ-<�}��tC<V�� ��<� f>��}=�<�~.�<2� .  P��X�~J�<�|��tC<V�� .� �|�=�<�~.�<2�.  ���XTJ-<�}��tC<V�� .> �}�=�<�~.�<2� .  ���X�}J�<�|<�tC<V�� ��<� f���|�=�<�~.�<2�.�  @ �X�}J�<�|<�tC<V�� .� �|�=�<�~.�<2�.�   � J�J�}9���~t=  `� ��f�~���J�t��<�	<�v �}t�<�~<C<�����t��<�	<�v �|�=�<�~.�<2�.�|<�< �~X Cf=�CX  P�v= JZ�X==$  ��.���}JN�<g�}<���}f���}X   �t� ��~<� <�<�z<� �/0MK�1K�J>�}</-=	.w�L�.==�}._  ��<�>�<�~<�.�{<��1�  ��<���� <�{X�<�{��  0� �j����zf�<�z<=�X�z<�J�J�|J/q�	� X��X�f�~t�K�.�<�<=;=��yJ2X�<���d=!e���~<�<C<�~�=�<�~.�<j	N���JV<*X����v<
t< 	:� 	Cf   ��J�~J�J�~.�;/�J�~<�.�{<u�  @� ��f�~9�~<�.�~.1>�<�~<�.�{<L�1<��CfV�   �t`� <
r<J`J
X�\.$J\<%</-Y�ge/j � t����}<�zX�i �\hH�f�}<v ��� et J�f= �}� x�z�=s�sKIuI2%  p	�t�<
<n�� X�t� <v �J n. �$���J�}< J?wvN��=�}�Z�X�}<g  �
���fK�~��<�}X���}<k<�t�~t�f��~�  p���<�I=�~��~<���}<k<�t�~t�f � _�  ����f�}<�<!�}��.�~f�~��<�}��<�}J�<�~��~<�<�~.2/H�f�~<�.�{<��d$CfV� �f�f  ����<�I=�|��<�~<���~t�<�}��<�}��<�~��~<�<�~. � 2< / H �f �~<�.�{<��d�CfV� � J4t  p�f�S��~<�tC<V��.���}�=�<�~.�<2  ��   ���f�~���J�t��<�	<�v �}t�<�~<C<� ��
��t��<�	<�v �|�=�<�~.�<2�.�|<�<�~XCf=�CX  ���X� J�J� .�~<�;/�J�~<�.�{<��  0��Zf� <�<'<*��}<k<�t�~t�f��}�   ��!<�I� fV<*��}<k<�t�~t�f � �~�   ��Hf:<F<:<.if�}��<�}��<�}J�<�~��~<�<�~.2/H�f�~<�.�{<���~$CfV� �f�f  `��<�I�}f�<i<�it<�}��<�}��<�~��~<�<�~. � 2< / H �f �~<�.�{<���~�CfV� � J�t  ��f��~��~<�tC<V��.���|�=�<�~.�<2  p�  ����~f�~���J�t��<�	<�v �}t�<�~<C<���	��t��<�	<�v �|�=�<�~.�<2�.�|<�<�~XCf=�CX  p��~X�J�~J�.�}<�;/�J�~<�.�{<��  ���� fK�~����}<�<�}��� ��<�}����~t�<�|"�f  ����<�I=�~�� X� <�<�}<���~t�<� �}�   ��6fK�~����}<�<�}��� ��<�~#�~<�<�~.1�O<3<,>�.�<�{<���|'��CfV� �J�|<��  ����<�I=�~�� X� <�<� t�<�~5�~<�<�~.1�O<3<,�<�~<�.�{<���|���CfV� �J �}���  ��f��|��t�}<DC<V��.�z<����|J=�<�~.�<2  0�  @���}f�~���J�t��<�	<�v �}t�<�~<C<���	��t��<�	<�v �|�=�<�~.�<2�.�|<�<�~XCf=�CX  0��}X�J�}J�.�|<�;/�J�~<�.�{<�� �   �  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  ios.cc   ios_base.h   atomicity.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   char_traits.h   c++config.h   cwchar   clocale   allocator.h   basic_string.h   basic_string.tcc   locale_classes.h   stringfwd.h   limits   postypes.h   functexcept.h   debug.h   predefined_ops.h   new_allocator.h   exception 	  locale.h   atomic_word.h   new 	  <built-in>      p�  M�8�|# J    �� ^Y%<[<&f   � J���}�  P � �Fi9@h�>V>�> ����}  J� � �� �gf*t;==g�wf<k<0g	tz<By�8h� �c<<c<)<W<1gwvf��w�   "��g=��z.R~y�	  p"�XK=�J=� <�.� <[;/c�t=� <�.� <4u  �"� J���� J�yt	twJ  0#� J	J |     �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext  locale_facets.cc   ios_base.h   basic_string.h   locale.h   clocale   cwchar   char_traits.h   stddef.h   c++config.h   allocator.h   basic_string.tcc   stringfwd.h   locale_facets.h   ctime   locale_facets_nonio.h   stl_iterator_base_types.h   stl_algobase.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   debug.h   predefined_ops.h   new_allocator.h 	  stl_iterator.h   cpp_type_traits.h   atomic_word.h   time.h   <built-in>      P#>X�hYuYm+=v/d�S`�g;1Y=*[=z�k=  �#� �<�~J�J�~.g�K� �ue�;ZvpJ ,   �  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  locale.cc   atomicity.h   basic_string.h   locale_classes.h   char_traits.h   locale.h   clocale   cstring   cstdlib   cwchar   cpp_type_traits.h   stddef.h   c++config.h   allocator.h   basic_string.tcc   stringfwd.h   ctime   stl_iterator_base_types.h   c++locale.h   string.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   functexcept.h   wchar.h   debug.h 	  predefined_ops.h   new_allocator.h   stl_iterator.h   concurrence.h   type_traits.h   gthr-default.h   atomic_word.h   time.h   new 
  <built-in>      p$�  �$�  �$� �  �$�   �$� �:>�.�~f����W�|t��t���z��.�}<�<=��y 2J�.���<�~<�t���z��.�<=��y 2J�.��� X�<� <���z��.�}<�<=��y 2J�.�t� <�<� ����y�	�� ����x�<X
t<YX
t<���x�
t<2�RC<�~=�<�~.�<2  @'� �l� ���Mw �� �~f �< �r. �<�nXC<=fC<=fC<�~�z 4 ��v<
X�����l =�<�~.�<2�~#=�<�~.�<j,1`C<�~�g�=�<�~.�<2  �(�<L JO� \�$tp�Y�Y�Y��  �)�>  �)��ut7X  �)�  �)��? ut f��~t=�<�}<�<2�~�� J� ut ���~t=�<�}<�<2�~�� J�� t Z J = s=��wB	  P+� Kjf/�<�|<�.�|.���|��J  �+� f�/V.y</�<�|<�.�|.0��|�0  �+��i�p@ = ; gJ���~� �J � � ; = - =���~� �Jz % �3��;=ua�}���  �-��;g� ��}f���.� <�f�9AV>�e/ � �L � s�@~@ m y< CJ � �� � s�9===+? .� t�}��<�}<�Jg�}f=�<�}<�<Y.`& zf��}J=�<�}<�<2g���4���� �	   0�X� ��}f���~.�<�~<u��WW  �0�<�  ; = ��  �0��}�t<�}��.� J m y<�}��J0�}�&  @1�K�}f��0= 	   �  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  streambuf   postypes.h   streambuf.tcc   char_traits.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   c++config.h   cwchar   clocale   allocator.h   basic_string.h   basic_string.tcc   locale_classes.h   stringfwd.h   ios_base.h   stl_algobase.h   debug.h   predefined_ops.h   new_allocator.h   exception   locale.h   atomic_word.h   new   <built-in>      `1�  p1�  �1��|J��  �1��|J��  �1�  �1�  �1�  �1�   2�  2�K  02�JK  `2� N*@F����|<t�kX���~X�.�~f�<�z<b�u�=m<   3�JN�w<	XyJg�~��~<�<�f  @3,N*@F����|<t���{�k����~X�.�~f�<�z<b�g�m<J�<�~<.�.g�~��~<�<  4��fq��=!  �4�KIK  �4� K  �4�X���� �5  P5�<��~���3  �5�"  �5� Lg g �     6�J�J?�~<�J�~fLJ<���|�7]'Y�'Jm�hf��g�~�  �6�J�J�~<bX�<�~fr�Ȝ�}�LH��g�~�  P7��J�~<LX7J"�  �7�K  �7� � ��<�'� ��~f� J�f� <�J� Jy   �7�<� J�<� X�~f� Jr  08� � ��<Z� .�~J�<d�~ �<�~f�J  �8�K  �8�M<  �8�  �8�  �8�   9�  9�Luu  09�  @9�  P9�  `9�  p9��g  �9�J�}J�<�}X�f�����~��JsKI  �9�   :�  :��=  `:�  p:�@! j     �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  locale_facets.h   basic_ios.h   basic_ios.tcc   ios_base.h   streambuf   atomicity.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   stl_iterator_base_types.h   char_traits.h   c++config.h   cwchar   clocale   allocator.h   basic_string.h   basic_string.tcc   locale_classes.h   stringfwd.h   streambuf_iterator.h   postypes.h   functexcept.h   locale_classes.tcc   debug.h   predefined_ops.h   new_allocator.h   exception   locale.h   atomic_word.h   new   <built-in>      ���  ���  �:�  �:�J  �:� K  �:� � ��   ;�  ;(<�x;=0� f�X  P;�Qzt	  p;�<�AZI  �;�  �;�  �;�  �;�  �;�  �;�HL=   <�  <�MI=>   <�  0<4JMI==�  `<�XL�� ��|<�Jg�|J=M����y"  �<�Xn��>7f�|<�Jg�|JJ>����y*  P=�gI��}<�J�|����K�|t�X��yJ  �=�YIK�|<�Jg�|�����|��X�y.  P>�JL=  �>�X����$�#w.:v]:�1�  p?� i9<�f�{����~<=� Jq���t�2   @� X�i�zJP7Luu==  p@�X>@e  �@>t�� � w =FP�� J�v�e= � կ�f�}J�<� fif�}<<><�<�}f�}<�<�{��� �$<=�~�\ =�=-���| ���|<���|f� ��|<��g�|J=�t�+��y- �   8  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  codecvt.cc   codecvt.h   locale_classes.h   locale.h   clocale   cwchar   char_traits.h   stddef.h   c++config.h   allocator.h   basic_string.h   basic_string.tcc   stringfwd.h   ctime   stl_iterator_base_types.h   c++locale.h   stl_algobase.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   debug.h   predefined_ops.h   new_allocator.h 	  stl_iterator.h   cpp_type_traits.h   atomic_word.h   time.h   new 
  <built-in>      @C;��  `C� �  pC� ��  �C�   �C�   �C� ��  �C�   �C1X>eg�f�~f�<�~<�f  0D1JL  PD%�.�}.�<�}J�J�}.�f�}f��f  �D+� �}.�<�}J�J�}.�f�}f�      �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  monetary_members.cc    locale_classes.h   locale_facets_nonio.h   locale.h   clocale   cwchar   char_traits.h   stddef.h   c++config.h   allocator.h   basic_string.h   basic_string.tcc   stringfwd.h   ctime   stl_iterator_base_types.h   c++locale.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   debug.h   predefined_ops.h   new_allocator.h   stl_iterator.h   cpp_type_traits.h   atomic_word.h   time.h   new 	  <built-in>      �D(  �D-XL�K
<v�K�uuuuuuuu=h � ��nf���t�yu  F� XL�K
<v�K�uuuuuuuu=h � ��nf���t�yu  @G� X=;g J�=e  �G� JK  �G� X=;g J�=e   H� JK �     �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include/sys /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext  fstream.tcc   fstream   basic_ios.h   codecvt.h   char_traits.h   streambuf   stl_algobase.h   postypes.h   istream   ostream   ios_base.h   stddef.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   types.h   file.h   wchar.h   exception_ptr.h   cwchar   c++config.h   cstdint   clocale   allocator.h   basic_string.h   basic_string.tcc   stringfwd.h   locale_classes.h   cstdio   basic_file.h   c++io.h   streambuf.tcc   basic_ios.tcc   functexcept.h   locale_classes.tcc   exception   debug.h 	  predefined_ops.h   new_allocator.h 
  locale.h   gthr-default.h   atomic_word.h   stdio.h   <built-in>    new   stl_pair.h      H�X�|���L�tq��I=@  �H�<O.fR�Jx<�~f�Js�v�h��1m�X�~f   I�A)P���  0I�f���f� f�J� <� ��~f� J���� �R #.d<�J�<�}��<�~t�J==�<*�h�4Xw��~fL:� .�.�J��===I;=�<=  �J�t�{<���� �k� f =�|���xV00=+iz
�H�r�}�k� <==,<�� t�}�:>� <==�<�.�~f�}�  �K�tO�r�ȆQ�~<����[<(��zgI/x f �\
��p<R.-4.z.=<uJX���Kk
�kV�- ZX��uDt;�d0a�.��<��~t�J==�}�Xe�� �K� <=�<g�X��~tSJ� <�~<�.�<��}t�J==�}�� ��f� .�<� <�<� t��](���=�<�}<�J�}<�<�}<���~f���~�� �D<�<��~t�J==�~<g� �s/i �==#� ���a<�K;Kt%�~�   P�yE�� X�}���<�}<�J�}<�<=� <K;=� � �{t����@�-K�/�s.��J�~�� J�J�<�� t�J==� <�<tJ.��~�� J�J�<�tEJ==� �1�<�}��</�}.�<�}.�X�~ȣ� J�J� <==,<!<t����JL:>� <==�<�.�~���D<?J9DX�}��J�}<�.0*�T�Z�|�   S�Lh?G=g�<=�}<  0S� Li���}<=H�f>�}<�<�}<  pS� ��<�}��<�}�s�W�� �  �T�
  �T.JO fy��I=  �T<JMh t�uL t�uuuu  @U��l�|<����	t�}<��=A��}f�X�}��<A�|.�t�|X�Ȅ
�.Y^�fu�t�$�|<���=;/�Yf��|�  �V�JM�{<�fuf�{f�<�{<��  �V��xY� � �y<�����z��� s� ���z<�<�zf�.0[g
Jz�]l�Yg�,XN���y�  @X�t�z����s��?Av.K�~J���|f�<�t�}<==�<
  �X�X�i�~f���I!��~X�fM�~J�J��=-g.:Xf�I���<�Qt==N<-K�~X�J�}��.�~.�Jh�~J���}.g�<�}<H�<>�}<����k� <==,<��~�:>� <==�<�.�~fU� <==,<�~f � �   �Z�t��|t����{�� J�<�{.���|��J�|.�X�|.�<Q �f�J��� ^t �{< ���{�ig�<�}<H�<>�}<���<��2k�e
J�y$B  �\�X�{��<� ����{J�f2�{�g�<�}<H�<>�}<��  �]�f��z���(J?X� � �y<�������y<������zJ��w�zf���u X�� ��{��<�Qt==����zf�<�zf�<�z<��73SAM=-=��x<  @_� �>h=� <=�<g\ ���t�~f?�t��~t� �  �_�  �_��}
  �_��}
  �_�   `��|
  `��|
   `�  0`��{
  @`��z
  P`�JL�Kg�.�}<K�J�Qt==�}<  �`� �� <���q<<t�>:uKg�<�}<K�J�Qt==�}<��;/V *.p���Zz ^  �a�JKj�<j��jJ  �a��	�f�~<	�<!�~�g�	 �}�  �b��<	�I=�~� t /t �~�  Pc��
�~f�<
�~<�<g�
 �{�  �c���~<
�I�f t /t �}�  �d��	�~fK
�~�	��h<	<h�	�z$�f �  �e���}<	�I=
�~��X�� � �{�  �f� f���~����������}<u�?K�JRt==,<u�|t	.e<.yfH��e<.  �g�  �g��|J�J�|J�<�t�}<�fyIT�|Xz<Pz<�J�|J  �g��{J�J�{J�<�t�|<�fyIT�{Xz<Pz<�J�{J  Ph�J�{J���{<�fyI��zXz<Pz<�J�zJ  �h��|J�J�|J�<OIp�|Xz<Pz<�J�|J  i��{J�J�{J�<OIp�{Xz<Pz<�J�{J  pi�JMyI��zXz<Pz<�J�zJ  �i��	�zfK
v�	��<	<�� 3�J� X�z.�<�zXzf�t�<	�z.�f �  k��	�zfK
v�	��<	q<��{��<�{<��O�J� <�z.�<�zXzf�t�<	�z.�f �  Pl���}<	�}I=
v��X�� �3�J�  �z.�<�zXzf�t�<F � �{�  �m���}<	�}I=
v��X��{t�<�{<��O�J� ��z.�<�zXzf�t�<F � �{�  o��
�}f�<
�}<�<h�{��<�{<�<�J� .�{.�<�{Xzf�t�<�
 �{�  �o��
�}f�<
�}<�<h�{��<�{<�<��O�J� �{.�<�{Xzf�t�<�
 �{�  �p��	�f�~<	�<!�~�h�}��<�}<�<�J� ��|.�<�|Xzf�t�<�	 �}�  �q��	� f�<	� <!��h�}��<�}<�<��O�J� X�|.�<�|Xzf�t�<�	 �}�  �r���~<
�I�f t 0�{t�<�{<�<�J� <�{.�<�{Xzf�t�<� �}�  �s���~<
�I�f t 0�{t�<�{<�<��O�J�  �{.�<�{Xzf�t�<� �|�  �t��r<	�I=�~� t 0�}t�<�}<�<�J� ��|.�<�|Xzf�t�<� �~�   v��b<	�I=�� t 0�}t�<�}<�<��O�J� ��|.�<�|Xzf�t�<� �~�   w�JL��|.�<�|<zf��  `w�JL��{.�<�{<zf��  �w�JL��y.�<�y<zf��  �w�JKjf   x�X��|�jt
� ��  �x�X��}�jt	� ��  �x�JK�|�jt� ��<� ����|J��  Py�JK�}�jt� ��<� ����~J��  �y�X��{��t�{fj	� 
�z<	���  Pz�JK�|�jt�  � �  �z�JK�}�jt�  � �  P{�JK�{fjt� ��<� ����{J�f�  �{�JK�{fjt�  � I� �$   N  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11 /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include  basic_string.h   stl_iterator.h   char_traits.h   basic_string.tcc   new_allocator.h   atomicity.h   stl_iterator_base_funcs.h   initializer_list   cpp_type_traits.h   stl_pair.h   stl_iterator_base_types.h   c++config.h   cwchar   cstdint   exception_ptr.h   allocator.h   clocale   stl_function.h   stl_algobase.h   functexcept.h   debug.h   predefined_ops.h   string-inst.cc   type_traits.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h 	  locale.h 	  atomic_word.h   new   <built-in>      p|�  �|�K  �|�
  �|���|J�J�|J  �|�oJoJ.�<�|.  �|��<�|J�J�|XOF   }��<�|֠I  0}���|J�J�}.�  P}�J6JJJ9.   p}���X`"  �}���Xd"  �}���X\�  0~�
JvJ
JR.�X`�  p~�JuJJM.�X`�  �~�KIKR.�X`�  �~�LHLM.�X`�  0��  @�  P��~  `��~J�  ��� �J� J�J  ���}�J�}J�.� <�.  ���}�J�}J�.�{<�.  ���{�J�{J�J  ��(XJ(JYJ  ���|�J�|J�.<a.  ���|�J�|J�.�{<�.  0���{�J�{J�J  @��
  P��
  `��  p��
  ����� f	  ����  ����{<�J�{J�.�<O/E  Ѐ�  ����z�f�<� J  ����|J�J�|��.�|<J�tK�}.�X��|f�f�|t  p�� �~��.�~t�.�}f� t�J�}�	  ���JM�  Ё�JL�  ���   ��  ��   ���|t�J�|J�.n.</�w�6xX 0�1K �|� �<%  ����s<�f  ��J�sJ���  @���|<�JU�|��.'<	J�|.�<�|.�<�|.���|.�<w  ����|t�J�|��.�X9<Jv���{���P73�Y   ���s<�f  @��J�rJ���  p���| �J�|X�.�X� <	Jy��K �]  ���
.vXX��{J�f� <�{��JGzY�1  0���r<�f  P��J�rJ���  ���  ����{t�J�{��.�.� <f;Yv���{�� P73   ���r<�f   ��J�qJ���  P��  `���{t�J�{��.�<�~.�J�{f� M:0�Y  І��q<�f  ���J�qJ���   ���{<�J�{��.�<��wY  p���{t�J�{��.�~X�<Jv���{�� P73�Y  ����q<�f  ��J�pJ���  @���{ �J�{X�.�~X�<Jv���yY  ����pX���}��~.���X  Ј��{<�J�{��.�|<JPt^J"<�.���|.�~.���X�{J  0���{t�J�{��.�|<bJ�f�|<J� ���zJ�����{�"  ����zt�J�zJ�.�|<� �~.���X   ���zt�J�z��.�|<J�t�.�{��~.���X�z�  p���zX�J�z��.�|<J�t���{.�~.���X�zf  Њ�  ���  ���   ��  ��   ��  0��M�vJ
t.  `��  p��J�#�4z< . � ="���|<���|<�t�X  ���OS<�N���~f?.�<�.�.T�� Y�
t.  p��>� ��f  ���>6.Kf  ���  ����}  Ќ��~J=�<�~.�<5��  �� Mt�~J=�<�~.�<5  @���~JnC<���|�=�<�~.�<2  ����~t���~J�.=<�}<=h��V0�~.� J�~<� <� .�~�J���~JnC<9�����t��X�����eK�J��_�z<
t<�J�~ $�~<=�<�~.�<j  P��J�~J�.wu�}�t  ����J� .u  ���X�}�.u���.
  ���X�}�.u�~��.
   ��X�}�.u��=� .�.  `��J�{J.u��K  ���J�{J.u��  ���X�{J�.�{fu���<� .  ��X�{��.�<�{Ju��;/z<  0��X�}�.u��<�{.�.  p��<K�.� .  ���
X�z��}Xn��J��w�  ���
<�|J�J�|J�.�w��.�vX�	t-/   ��J
JvJ
JR/���|���� f�J�{<�tN  ���t:<�|����u�}.�X�.�|t�J�}�  ��	=WK�|X�.  @���J�{X�J�| �.�{�  p��
J��{X�|X�J�xX  ���
<�|��J�|<�.�w�.�vX�	t-/   ��t��yX�}Xn��	J�v�  `��T��zJ�f�zJ�.	  ���	�<�|X�J�zt�f�|t  ���<��u�}.�X��|��.  ��<#�(.�f�|<f��sJyK� J�X��z�
t<�� J�Xd�� f  Е�JL�  ���y<�J�y��.�}<n��J�yX  @��J�yJ���  p��	  ���J�}J���{�  ���t���.�|<
��J\�fz;/-/�X� .:=/pt�X� �v�NjJ���.h���� ������~<�.�f1S
  0��	�}J�f	  P��	�xt�J�x��.�}<n��J�x�  ���
J�wJ���  ���	�x<�fg   ��<�zJ�X�w<�J,��wJ  @��MZt*<�~.�J*<  `��<P�hgWY�}J�~<�<�~.4<� ���|<!fl<sJz.
t.�X  ��t�~��.�X�~<�~��<�~�K.=<C<9��.v��|�=�<�~.�<j  ���f�|<�.���+�  К�ta��.�|<]J�.�|<=Y=.�X��.� tz��.Y�
t<  p��  ���Pt0JP��.�|<�yKJ�.�}<=YuQ�X��.�tz��.Y�
t<� f  P��t�xJ(.�X�|<c�=-XVJ(*.��2.�.� tq -t��� �Zf;/mtX��
t<� f   ��  0��J�zJ���  `��  p��J�zJ����  ���t�
J(.�X�|<Qf=Y!� .�X.�.� tz�T�Y�
t<� f  P��J� ��|.�X�|<�.L1�}��.�z��F�}X  О�=  ��<�y��.�<=��y 2X�.�t�y
t<�J  `��<�z��.�<=��y 2X�.�t�z
t<�J  П�^�%< JZtCs�~�   ��� <�f� <�< J��f7�..�f�t  ���f3JP�KJ� <�< J(�C<9�U.�~�=�<�~.�<2l.�~�  ��   ����|���fg.��|�CX  �����|��fu.�-=נ�|�CX  ���?���o�CX  `�� t�
J�<�y.�f�y.�f�~f� .�<�.��B�� ���m<X8�
t.  �� t� N�OV<*.Vf*.�f�~f� .�<�.��B�� ���m<X8�
t.  ���� X�J� ��.�}<�~��J�J�s.�.�t��f�f  ��J�t��|X�J�qJ  0��� X�J� ��.�}<�~�� J�J�.�t��f� f  ��� t� N�OV<*.Vf*.�f�~f� .�<�.��B�� ���m<X8�
t.  0��<�J�tf�f�tt�f  `����� <�f�.�|<�x��� �<n<v�W��~��<�~<C<�~�=�<�~.�<\����~��<�<�<�.�J���X�~�t��tv� i. Cf   ���v<�	f  0���vt�	J�v��.�}<n��J�w"  ���J�vJ�	fK  Ч��zJ�J�zJ�.�zJ�.	  ���v<�	J�v��
.�zJ�f�z �.jt   ��<�u��
��zJ�f�z �.t=  `����zJ�J�zJ�.�zJ�.	  �����zJ�J�zJ�.�zJ�.	  ����yJ�J�yJ�.�zJ�.	  ����zJ�J�zJ�.�zJ�.	  ����yJ�J�yJ�.�yJ�.	  @��#U<M0JP� �. �t� Ef  ���<�J�sf�f�ttZf  ���  ���  Щ��<�t.Sf  ���<�t.Sf  ���<�t.Sf �	   �  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11 /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug  basic_string.h   atomicity.h   functexcept.cc   exception   new   typeinfo   system_error   future   functional   stdarg.h   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   cstdlib   exception_ptr.h   c++config.h 	  cwchar   char_traits.h   cstdint   stl_pair.h   allocator.h   clocale   basic_string.tcc   stringfwd.h   initializer_list   uses_allocator.h   tuple   ctime   chrono   mutex   shared_ptr_base.h   regex_error.h   stl_iterator_base_types.h   debug.h 
  predefined_ops.h   new_allocator.h   stl_iterator.h   concurrence.h   wchar.h   locale.h   atomic_word.h 	  time.h   <built-in>      0���~J=�<�~.�<5U  `�6<�kf  ��:<�h  ��><� ��f  �� <���~f   �� � �" �~< �< C<�~t ��.Cf  ��� � �" �~< �< C<�~t ��.Cf  @�� � �" �~< �< C<�~t ��.Cf  Ь� � �" �~< �< C<�~t ��.Cf  `�� � �" �~< �< C<�~t ��.Cf  �� �=igT@[9N*@u �( �~< �< C<�~t ��.Cf  ��� � �" �~< �< C<�~t ��.Cf  @�� � �" �~< �< C<�~t ��.Cf  Я� � �" �~< �< C<�t ��.Cf  `�� � �" �~< �< C<�t ��.Cf  �� ��"C<=<C<�t0  `�� �=�"t��n�<n<C<�t�<�~����~<�$Cf   ��`f <<O�t���~<�<C<�t`< �`� f �.Cf  ���<	���sf  в�X= <   �  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include  regex.cc   basic_string.h   atomicity.h   exception_ptr.h   cwchar   c++config.h   char_traits.h   cstdint   allocator.h   clocale   basic_string.tcc   regex_error.h   stl_pair.h   exception   debug.h   predefined_ops.h   new_allocator.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h 	  locale.h 	  atomic_word.h   new   <built-in>       �#  0�#J  `�Ye<=�J�}<�<C<�~��!�=�<�~.�<2, `C<�~=�<�~.�<2    �  �      ../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include/sys /opt/MeetiXOSProject/MXlibraries/include  compatibility.cc   streambuf   char_traits.h   basic_ios.h   ios_base.h   c++config.h   cwchar   clocale   istream.tcc   istream   cstdio   postypes.h   basic_ios.tcc   debug.h   predefined_ops.h   new_allocator.h   cpp_type_traits.h   stddef.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   types.h 	  file.h 
  wchar.h 
  locale.h 
  stdio.h 
  stl_algobase.h   <built-in>      �<�=�=;u��z<l��L�f�~�xs����z.�X�.�z<�<Lf�~< ��<vXIt5�*fV<%XOU��o�g�Xfc<#Xzff�`��f�~.�<�.�~fLt7X�}f?���h��,��~��.fR<)XOgO �.XTt �    �   �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  bad_cast.cc   <built-in>    typeinfo     p�  ��  ��J K   _  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits  vmi_class_type_info.cc   cxxabi.h   tinfo.h   typeinfo   stddef.h   c++config.h   <built-in>      ��K  жJK�   �$tKIK1��X�}X �xJ<b.fn./n�XY 7XJ���� XCJi�  �� tKg� ���v��VWU�w�7#��� .�~�#X]�#J�J�}X8NK.6JJJ.-.GJ9JLY�Z�B�HsL=W;Yf�	��9?ul��!X�	�-=hW��MJh� ��u�A<���� JKgV=y%E<s�KL+=>�l.� ���� J�J��� J4�J���� J<��~ � � KJ���i�LH=K-=f.��.�~�H�,u���T�~<�t�~<�.�~�L�=�ta�uuj�qtDt<X�X6��A�96Df  `��u"u-Ki(�  �}<xJft.�J��u�~X�Juv���L�~��#*2*G<2��;�1L+<q�K�~����cLY�� �c��t
 y    c   �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++  del_opv.cc   <built-in>    new     ��    �  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  eh_globals.cc   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   cstdlib   exception   unwind-cxx.h   unwind.h   <built-in>    cxxabi.h     ���  ��� �   �  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  eh_catch.cc   unwind-cxx.h   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   cstdlib   exception   unwind.h   cxxabi.h   <built-in>      ��u   �(<M�X�~X�~<�.�}��N2.h�?192=LL=�.�}<l.r�  ��� KY2�J�~ Zf�CeX_=Q_\=qtY�z   ��=Y� �     �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits  eh_exception.cc   cxxabi.h   cxxabi_forced.h   exception   <built-in>       �  0�  @�&  P�/  `�  p�  ��   ��   ��"  ��" 6   �   �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  tinfo.cc   typeinfo   tinfo.h   <built-in>    cxxabi.h     ��  ��8  ��?  ���    �  �� 4��NX2 NX    �   �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include  class_type_info.cc   tinfo.h   typeinfo   cxxabi.h   stddef.h   <built-in>      `�/J� ���:�HJ-9<G<ZYY  ��>!  ��K  ��JK�   �� ��pJ.Y�qJz�KvWr4  ��#t� X���J,\E]�s  �� XKIu,���cJ �JY�].KI/=xu��'X �    e   �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++  bad_alloc.cc   <built-in>    new     ��  ��  ��J V   �  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include  eh_terminate.cc   exception_ptr.h   cstdlib   cstddef   c++config.h   exception   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   unwind.h   <built-in>    unwind-cxx.h   cxxabi.h     �+[KZ��y.	  P�7$<]X  `�==K  p�� 2<OX  ��� �  ��� ^  ��� �  ��� ^ 7   �  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext  guard.cc   cxxabi.h   exception_ptr.h   <built-in>    c++config.h   cxxabi_tweaks.h   exception   concurrence.h     ���<tJ[jfJ� X�X� .�J���|f  ���~	   ���~J�J b   �  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext  eh_alloc.cc   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   cstdlib   cstring   exception   c++config.h   string.h   unwind.h   unwind-cxx.h   gthr-default.h   <built-in>    concurrence.h   malloc.h   cxxabi.h     0�� [uhV0.�;=kJcihM;/
Xz�u;�  ���N�iU?�  ���NvV0.�jg-1M;/
Xz��  `��N��U?w	 �   �  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  new_op.cc   new   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   cstdlib   exception_ptr.h   c++config.h   exception   malloc.h   <built-in>      ��*%S<O2YL/y<g
tzX�c �    �   �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  bad_typeid.cc   <built-in>    typeinfo      �  0�  @�J �    �   �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  guard_error.cc   <built-in>    cxxabi.h   exception     p�  ��J �   �  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include/sys /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/MXlibraries/include  pure.cc   unwind-cxx.h   stddef.h   unwind.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   types.h   <built-in>    cxxabi.h   exception   unistd.h     ��/=�  ��6=� y   �   �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  dyncast.cc   tinfo.h   stddef.h   <built-in>    cxxabi.h     ��0t�uJK.l<� <��.� .���.JRX[+�U<5XO<]sJ.� ��J� .�JM�  Z�.
 ;   �  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include  eh_aux_runtime.cc   typeinfo   new   exception_ptr.h   cstdlib   cstddef   exception   c++config.h   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   unwind.h   <built-in>    unwind-cxx.h   cxxabi.h     ��!<���~f  �%<���~f  @�)<�cf  p�-<*�Vf �     �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include  si_class_type_info.cc   typeinfo   tinfo.h   cxxabi.h   stddef.h   <built-in>      ��K  ��JK�  ��2t� 6=�DȦ8sp�I/=�nJ�s�u ?�J��H�u   �$t=L�s � <J����  ��� t���us 
     �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  unwind-cxx.h   unwind.h   exception   <built-in>    eh_term_handler.cc   cxxabi.h    �   D  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/MXlibraries/include/sys  vterminate.cc   typeinfo   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   cstdlib   cstdio   cxxabi.h   types.h   file.h   stdio.h   <built-in>    exception   malloc.h     �,��xY+�ZX&t]X؎0ד>�uXl.=�5���/���XVu�� &   �   �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include  eh_type.cc   unwind-cxx.h   cxxabi.h   unwind.h   exception   <built-in>      ��$=Y/Ll2z��.�~� 
     �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  unwind-cxx.h   unwind.h   exception   <built-in>    eh_unex_handler.cc   cxxabi.h    �   ]  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits  bad_array_length.cc   exception_ptr.h   new   <built-in>    c++config.h     ��   ��  ��J ?   �  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  locale_init.cc   locale_classes.h   locale_facets.h   locale_facets_nonio.h   atomicity.h   basic_string.h   locale.h   clocale   cstring   cstdlib   cwchar   char_traits.h   stddef.h   c++config.h   allocator.h   basic_string.tcc   stringfwd.h   ctime   stl_iterator_base_types.h   codecvt.h   c++locale.h   string.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   wchar.h   debug.h 	  predefined_ops.h   new_allocator.h   stl_iterator.h   concurrence.h   cpp_type_traits.h   gthr-default.h   atomic_word.h   time.h   new 
  <built-in>       �!>�  P��&z�M9?�+vu v �\u�v���
X�. � �~.��< � �. �ut �	� �vb �
� =X�w< � �~< �� �u���~<���r��~.��P�0<PX�~.��� ����{���=�|� � �~< �� � � �� �{� �� =X�|< � �~< �� �y���~<�	��x��~.�~����}����� � �~< � ����~<���~��~ �� �� Y Y Y � y< {�J�}����z��{�	  0��?Y�  `��7Y�  ���  ���J� �G�u�~����~X�<0�~f�<   ��<m��"  `��,�Tf,<�~���;id�~.�<-g�X�n�2JDC<��w�1�nC<�~�=�<�~.�<2,�`C<�~=�<�~.�<2    �  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug  ios_failure.cc   basic_string.h   atomicity.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   char_traits.h   c++config.h   cwchar   clocale   allocator.h   basic_string.tcc   stringfwd.h   ios_base.h   exception   debug.h 	  predefined_ops.h   new_allocator.h   locale.h   atomic_word.h   new   <built-in>      ��*  ��%X�J�~<�fC<�~���=�<�~.�<2  ��%JK   �"�=;	 �   �  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext  ctype_configure_char.cc    locale_classes.h   locale.h   clocale   cwchar   char_traits.h   stddef.h   c++config.h   allocator.h   basic_string.h   basic_string.tcc   stringfwd.h   ctype_base.h   ctime   stl_iterator_base_types.h   cstdlib   cstring   c++locale.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   debug.h   predefined_ops.h   new_allocator.h   stl_iterator.h   cpp_type_traits.h   atomic_word.h   time.h   stdlib.h   string.h   ctype.h   <built-in>      P�*  `�,� �}f���}X8�.�}<:@8N:�,vb@v�K$u   �8� �}f���}X8�.�}<:@8N:�,vb@v�K$u  ��� <  ��� X�0g;�P  �� <  0�� X�0g;�P 8     �      /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext  collate_members.cc    locale.h   clocale   cwchar   stddef.h   c++config.h   ctime   cstring   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   debug.h   predefined_ops.h   new_allocator.h   cpp_type_traits.h   time.h   string.h   <built-in>      ��+=ɟ;/  ��4 �   �  �      /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include/sys /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  stddef.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   types.h   file.h   wchar.h   c++config.h   cwchar   clocale   cstdio   globals_io.cc   debug.h   predefined_ops.h 	  new_allocator.h 
  exception   locale.h   stdio.h   <built-in>     �      �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  istream   basic_ios.h   iomanip   ostream   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   cwchar   clocale   char_traits.h   c++config.h   basic_ios.tcc   locale.h   debug.h   predefined_ops.h   new_allocator.h   atomicity.h   new   <built-in>      ����{J���   ��J�{J��t�  P��K	  `����z�Kv����z.�< �z�  �����}f�}F=v� �J �z� �< �{  ��� �z����   ��X�~f;K�~����|.�< �zt  �����}<�F=�~� �X �|� �< �{ �     �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  numeric_members.cc    locale_classes.h   locale_facets.h   locale.h   clocale   cwchar   char_traits.h   stddef.h   c++config.h   allocator.h   basic_string.h   basic_string.tcc   stringfwd.h   ctime   stl_iterator_base_types.h   c++locale.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   debug.h   predefined_ops.h   new_allocator.h   stl_iterator.h   cpp_type_traits.h   atomic_word.h   time.h   new 	  <built-in>      P�'XL�uuLK� � �� x ���uuumf���	t�s@  P�� X=;g J�=e  ��� JK �   �  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  locale_facets.h   istream   basic_ios.h   istream.tcc   ios_base.h   streambuf   char_traits.h   ctype_inline.h   postypes.h   iomanip   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   c++config.h   cwchar   clocale   allocator.h   basic_string.h   basic_string.tcc   locale_classes.h   stringfwd.h   ctype_base.h   ostream.tcc   basic_ios.tcc   stl_iterator_base_types.h   streambuf_iterator.h   stl_algobase.h   functexcept.h   locale_classes.tcc   debug.h   predefined_ops.h   new_allocator.h   type_traits.h   exception   locale.h   atomic_word.h   atomicity.h   <built-in>    new   ctype.h     ���  ��� K���~�   �� J�J�~<���~��  P��  ��Iu  ��� ��<�}@=�t   �� �  @��   P�� JL�  p��JL�  ���  ���XK.�|t�J�|����y%   �� �=  `����~<�@=�}f  ��-t�?0K��� �Pz.�J� t�X ����}��<�~<.t< f�X���~fL� �~<��J!zy��<�~.q��KM�!tY�!XzbXtqtt91\ $t�<h�+'�}��f�} ttttX  ��� k7<A��*x�����q*�<�q<tg<�g<%<l<Nmtl<�l<<.l<//;_z<�s���� ��.n<<OgpX�.r<	XOqf�XkX�  @��k7<A��*x���t�q*�f�q<	.xqT.,<ZXz</��~����e.<`<OgX�a.<\XOf�eXX�  p��\8<j�����.� <�Xz<� ��x#�G.9<B<Og;X�C.=<�XO<f�GX6X�  ���Qy<<Av��� �bX�<�~ftxX��.� <�XO� �1��.� <�<z<� �:����x֒�.� <�<Og� ��X� X�  ���O7<?v����~.�<�~Xz<��it&�bX�<�~f>r*�V�Xx.��~.�<�~<Og�X��~.�<�~XO�f��~X� X�  �����:v�g����k��T<-�wJ�J�~fLJ"<�~���u=�~t�<�~.�<�~Xz<��f�h�W�$�Mo���~.�<�~<Og�X��~.�<�~XO�feX��~X�X�  ���XK� .�|t�J�|����y%  ��k7<iv���� �f�L�� <����� .�~�HJ���~f.RXӑ�~.�<�~XO�����~.�<�~Xz<����h�+<� 0�~f�<A�e��e<.���~.�<�~<Og���~X�X�   ��XK8.�|t�J�|����y%  ���N8<?u��n��~��Xift�~ ��X�}.�<�}Xzf���}.�<�}<Og�X��}.�<�}XO�f��}X�X�  ���O7<@u���}�LX�<�}f��X�|.�f�|<zf��zX��|.�<�|<O�fo���|.�<�|<Og���|X�X�  ���N8<?u��q��}.��;=.�{.�<�{Xzf�t�{.�<u���|.�<�|<Og�X��|.�<�|XO�f��|X�X�  ���N8<?u���|�g�JK�}.���}<�<r���|���<�{.�<�{Xzf�<��{.�<�{<Og�X��{.�<�{XO�f��{X�X�  ����m,v�{X�fu喟�}t��.� .�<� <���{�z<Bz<���~��Ȓ�{.�<�{<Og�X��{.�<�{XO�f��{X�X�   ��tC,v�{X�fu喟�}t� X�f�}t���{ z<Bz<�t�{.�<u���{.�<�{<Og�X��{.�<�{XO�f��{X�X�   ��Pz<<B����{J��[.eX��z.�<�z<zf��Xu���{.�<�z<Og�X��z.�<�z<O�fkX��{X�X�   ��^z<<	�zf�ȑ���{X�J�{<�<�w��z.�<�z<Og�X��z.�<�z<O�f��zX�X�   ���B�zt�fu���{���{f�<X�z.�<�zXzf���z.�<�z<Og�X��z.�<�zXO�f��zX�X�  @�����zt�fu���zt�<�zf�<X�z.�<�zXzf���z.�<�z<Og�X��z.�<�zXO�f��zX�X�  `��  p���}f�<C�}���0�zf�<�z�L� �~< w����Q�z����~��}��<�~<J�<�~.q�KM�!�Y�!��b��qt�q1\�$��th����yf�<�yXzf�t�y<�<�z����z<�� �  � �O7<A��o�{�bX�<�~f�X�{��X�y.�<�yXzf���y.�<�y<Og�X��y.�<�yXO�f��yX�X�  ��  ��   �  � 
  �<L�tf
�~��<�|<�J�|fnXJ
�~<�t��y� 
 �� Li�
t 
 �� LX
qJ.t.
; 
 �� � X � � Ft j
 ;X 
 0��J
�|J�.
�|t 
 P��J
�|J�.
�|t  p� i9<?��+wQ��J�q,x..R<4Xz<U�D�1��?.A<:<OgCX�;.E<6XODf�?X�X�  ��  �� i9<?��+wQ��J�q,x..R<4Xz<U�D�1��?.A<:<OgCX�;.E<6XODf�?X�X�  ��  �� i9<?��+wQ��J�q,x..R<4Xz<U�D�1��?.A<:<OgCX�;.E<6XODf�?X�X�  ��   � i9<?��+wQ��J�q,x..R<4Xz<U�D�1��?.A<:<OgCX�;.E<6XODf�?X�X�   �  0� i9<?��+wQ��J�q,x..R<4Xz<U�D�1��?.A<:<OgCX�;.E<6XODf�?X�X�  P	�  `	� i9<?��+wQ��J�q,x..R<4Xz<U�D�1��?.A<:<OgCX�;.E<6XODf�?X�X�  �
�  �
� i9<?��+wQ��J�p,x..R<4Xz<U�D�1��?.A<:<OgCX�;.E<6XODf�?X�X�  ��  �� i9<?��+wQ��J�p,x..R<4Xz<U�D�1��?.A<:<OgCX�;.E<6XODf�?X�X�  ��  �� i9<?��+wQ��J�p,x..R<4Xz<U�D�1��?.A<:<OgCX�;.E<6XODf�?X�X�  �   � i9<?��+wQ��J�p,x..R<4Xz<U�D�1��?.A<:<OgCX�;.E<6XODf�?X�X�  @�  P� i9<?��+wQ��J�p,x..R<4Xz<U�D�1��?.A<:<OgCX�;.E<6XODf�?X�X�  p� ?     �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  ios_locale.cc   stddef.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   char_traits.h   c++config.h   cwchar   clocale   allocator.h   basic_string.h   basic_string.tcc   locale_classes.h   stringfwd.h   ios_base.h   ctime   stl_iterator_base_types.h   debug.h   predefined_ops.h   new_allocator.h 	  stl_iterator.h   exception 
  locale.h   atomic_word.h   time.h   <built-in>      �&XOGuv;ug  �1<�ɻ�= �   �  �      /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include/sys /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  basic_file.cc    stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   types.h   file.h   stdio.h   cstdio   cwchar   postypes.h   c++config.h   clocale   ios_base.h   basic_file.h   c++io.h   limits   gthr-default.h   wchar.h   debug.h   predefined_ops.h   new_allocator.h 	  exception 
  locale.h   fcntl.h   time.h   stat.h   unistd.h   <built-in>    errno.h     � /-lzt<�Mv.� ��KW/  p�K  ��<������~�y/kp�.  ���~t�<�~<� �. wJN;KK�st	  ���~J�J�~J� �q<.x<[O  ��  ��f�	   �  0�XtJ.Ml�Ǐxk73}kl<.  ��  ��Np<$�;�  �X  @�/-<ON�91z��,02  ��Xm�vJ	   �  �X!J/@*K# �   �  �      /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext  messages_members.cc    locale.h   clocale   cwchar   char_traits.h   stddef.h   c++config.h   allocator.h   basic_string.h   basic_string.tcc   stringfwd.h   ctime   locale_facets_nonio.h   stl_iterator_base_types.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   debug.h   predefined_ops.h   new_allocator.h   stl_iterator.h   cpp_type_traits.h   atomic_word.h   time.h   <built-in>      `(J �   �  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include  stdexcept.cc   basic_string.h   atomicity.h   char_traits.h   c++config.h   allocator.h   cwchar   clocale   basic_string.tcc   stdexcept   stringfwd.h   exception   debug.h   predefined_ops.h   new_allocator.h   cpp_type_traits.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h 	  locale.h 	  atomic_word.h   new   <built-in>      �*  ��   �&X�J�~<�fC<�~�.=�<�~.�<2  �/   /J  04  @4J  p9  �9J  �>  �>J  �&J  � X�J�~<�fC<�~�-=�<�~.�<2  `�   p� J  ��   �� J  ��   �� J   � J  @#X=2  �,JK  �1JK  �6JK  �;JK   � X=2  @� JK  `� JK  �� JK �   �  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/MXlibraries/include/sys /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  c++locale.cc    cstdlib   cstring   cstdio   clocale   cwchar   char_traits.h   c++config.h   allocator.h   basic_string.h   basic_string.tcc   locale_classes.h   stringfwd.h   ios_base.h   ctime   stl_iterator_base_types.h   limits   c++locale.h   functexcept.h   debug.h   predefined_ops.h   new_allocator.h   stl_iterator.h   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   stdlib.h   string.h   types.h 	  file.h   stdio.h   locale.h   wchar.h   cpp_type_traits.h   atomic_word.h   time.h   new 
  <built-in>      �2��;/�Ƀ	� � ���%��p� �	��H�	  �� ��;/�Ƀ�82 �"u'��r� ����-]�	  ���hH�Y;/�׃��/۟�r�;K��gs sX��Vt	  �2�?KIgMe  P�  `�  p� �   5  �      /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++  time_members.cc    locale_classes.h   locale_facets_nonio.h   locale.h   clocale   cwchar   char_traits.h   stddef.h   c++config.h   allocator.h   basic_string.h   basic_string.tcc   stringfwd.h   ctime   stl_iterator_base_types.h   cstdlib   cstring   c++locale.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   debug.h   predefined_ops.h   new_allocator.h   stl_iterator.h   cpp_type_traits.h   atomic_word.h   time.h   stdlib.h   string.h   new 	  <built-in>      �,�=�;/�׃�   K � �u=qX	   =JL�uuuuuuuuwuuuuuuwuuuuuuwuuuuuuu�����������������G���~t�� �   d  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include  functional.cc   functional   exception_ptr.h   cwchar   c++config.h   cstdint   clocale   stl_pair.h   uses_allocator.h   tuple   exception   debug.h   predefined_ops.h   new_allocator.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h 	  locale.h 	  <built-in>    new     p!"  �!�  �!�J    l  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11 /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug  snprintf_lite.cc   stdarg.h   cwchar   clocale   c++config.h   cstdint   exception_ptr.h   ios_base.h   functexcept.h   locale_facets.tcc   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   locale.h   atomicity.h   debug.h 	  predefined_ops.h   new_allocator.h   <built-in>    stl_pair.h     �!1%S]�f>?4wf5yfCy<m0VM9>��  @"� $*NBwq?e/1!=F  �"� wMH2*tV� t�g�Nh ���{k<<tX1�=ggf��Kuu3y<R
� o   �  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/MXlibraries/include  future.cc   system_error   basic_string.h   atomicity.h   exception_ptr.h   new   stl_pair.h   cwchar   c++config.h   char_traits.h   cstdint   allocator.h   clocale   basic_string.tcc   stringfwd.h   initializer_list   uses_allocator.h   tuple   ctime   chrono   mutex   shared_ptr_base.h   stl_iterator_base_types.h   future   exception   debug.h   predefined_ops.h   new_allocator.h   stl_iterator.h   atomic_base.h   concurrence.h   stddef.h   stdint.h 	  fs.h 	  kernel.h 	  ipc.h 	  kernquery.h 	  wchar.h 
  locale.h 
  atomic_word.h   time.h 
  <built-in>      �#  �#  �#J  $�    $� J  P$� �� ���<�~t���w��X�y.�<�y<C<�~�=�<�~.�<2�����~<�<C<�~����yX`C<�~=�<�~.�<2  �%"�i�<�~f� �w.�.�w.m��X�w.�t�w.���w.��RC<�~=�<�~.�<2  �&� v
�v�
8	 �   G  �      ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11 /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/MXlibraries/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/debug /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/ext  system_error.cc   system_error   cstring   cwchar   exception_ptr.h   stddef.h   c++config.h   char_traits.h   cstdint   allocator.h   clocale   basic_string.h   basic_string.tcc   stringfwd.h   initializer_list   stl_iterator_base_types.h   string.h   stdint.h   fs.h   kernel.h   ipc.h   kernquery.h   wchar.h   exception   debug.h 	  predefined_ops.h   new_allocator.h 
  stl_iterator.h   locale.h   atomic_word.h   new   <built-in>    stl_pair.h     @'%  P'4  `'� � J��  �'�  � 
  �'1  �'"  �'1  �'"  �'8JNu	   ()JNu	  P(�  `(�J  �(� X� ��J���~t�J�~.���~�  �(�    )�   )�    )�   0)� J� ��X'  ��� \<=#f E     �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits  new_handler.cc   exception_ptr.h   c++config.h   new   <built-in>      �).�  �)=^ �   Z  �      ../../../../gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/bits /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/libsupc++ /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/include/i686-mx/bits  bad_array_new.cc   exception_ptr.h   new   <built-in>    c++config.h     �)   �)  �)J +   �  �      /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/../include /opt/MeetiXOSProject/temp/gcc-4.9.1/libstdc++-v3/../libiberty /opt/MeetiXOSProject/MXlibraries/include  cp-demangle.c    stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   demangle.h   cp-demangle.h   string.h   malloc.h   stdio.h     �)�zXl8J�J)<W.Zge� JNH/=[��+JV�?�.��~<�ge�<"g=�Xr0��f374-=  �J[Gl�-/>>`f�KL[G�L[G,.c .iȄ��tp<L�|p<./v�u�.282=�pXRI],>,>�sI���� . �f M 9 ? ?f).��=�v ��l��. �� ��	<w.uyM � �Vw.����?�L/f��7J�i��f�i<s�.�iJ0ge�<MIh;=�thL=C�i<�ge�<�g=� = �X�X-t/[� ��<� J�=�ȃ=f�=�fg��K�gq�;u�V��mf6x.Q/-=
X91l=WLxJ
�o<=�/ �y���y ge�<L���y�.�y��.�	�":0vwZ~_w� 4 i)f�	. sf # 9 # [ YM�oJ�ge�<M;g�.�q<�.���^7�Y+�q<\Y-/=f>�Ek5Yf��>� .Y�Y��Y��?���-.//�4 n֒Z�u � > , >zXX����>,c<NZHZFBx<
f�.m��~J�� �M.�L\<�.`u JX�|�<q�;KMts�//;�<L�zKW�-M�	t/q�{�gv;u�X�y�t��	�x.nt.fs<vf�+uht��y�y�t�Xw<	�x.nt.fsXv��,uh$"���t.fk��J;/�g&.��v�?�	��v<�	t�v�?�	��v<�	t��� <�w��<;hW�)AY J��{fBx<NZ�1�<�K�zt�
�v�!����xX!����X=-��w���;9�Ju�f=�gY�v*�	�xfntffs<v.uh�f���X���u#�	�xfntfXs<v.uh4�	�xfntfXs<v.uh4�	�xfntfXs<v.uh4�	�xfntfXs<v.uh"fy�ytCyXt�Xw<	�x.ngs<XsJv.uh4�	�xfntfXs<v.uh�	f�vf?��	�!��~Xgi*@���N ��x��	�xfntfXs<v.uh�f��x�	�xfntfXs<v.uh4�	�xfntfXs<v.uh�f����x+�	�xfntffs<v."Uuh� g>K����OX�矼��x*�	�xfntfXs<v.uhof����p�0��ۻ;/��.>1�ɻ
t��;AT=:>=9?>
 ������~�h@9q==;ih:>xu���9j=r�jx.>>@g>V�V\v�N8���xl.t\:h��W=�B��� ��W���~X��yX��yX��yX��yX��wX�!��wX��yX��yX��zX��X��uȅ	�xfntfXs<v.uh��� ��iH��h�XfEgx�=Bz<	f>/g��ʻ�ʽ���X�{�tȅ	�x.ntfXs<v.uh(�	�xfntfXs<v.uh�f!��g��aXK;g�}ft<�	�x.ntfXs<v.uh�fg�?g�83>zXg>;{=�j<v�|���Ldg�zXt��	�x.ntfXs<v.uh�f�}<�.=(����;?rgh�h��>,hg�~ֻ�yX��yX��yX���}��t0vZ:\ x��}f�}ȅ	�xfntfXs<v.uh�f���zX�䟻�-<�zX��}�N�x�t�	�x.ntfXs<v.uh�f�zX��X�v�?��	��� tɻɻ�zt�{)�	�xfnt.Xs<v.uh�f�\�\���;g� ���~�� =-=�vJ�	�xfnt.Xs<v.uh"fyfy4tXXw<	�x.n/s<XsJv.uhnٟ~�	�xfntfXs<v.uh�f��zftX�	�x.ntfXs<v.uh��=����y֯�.�	�xfnt.Xs<v.uh��=�37A*N���yX_ ��wJ�<�w<�f�w<�J�w.�t�wX��tu$Xt�la�;?x9�>g/r. ���|.�.Y�z����x<�t�x.�t�wX�r��K0,g�� ��~X�|�Bx<��\i�<�~��<Y�ut?��
f�/;uYglODs<Js.�ػ�uXuho������}��u�Vuh��u�V�u��Xh@9q==@7ih:>w���� ��g;��T�T�T�X��|.<iq=A)gh��.��y�z�����o���!���wX�u�����=�T�%>k98kolz<	�n<T�ʕ�-=L��XO���/�z>:=)������Hh���w �uh��w���w��wX�uh��uh�廻����x<�uh��uh�	��{X�}.�t�x��|���!��X^��X�uJ�
��u.u.u0s�<�;��	�"���u�t�?���t.�t-Xq�s��	�xfntfXs<vf;u"�#�t�	�xfntfXs<vf;u"3�	�xfntfXs<vf;u"3�	�xfntfXs<vf;u"#M�pٟ� �s�M���	�xfnt.Xs<vf;u"�'�t�?�I�	�xfntfXs<vf;u"3�	�xfntfXs<vf;u"�#�t�?��t�t"�	�xfntfXs<vf;u"�#�s�?�rX;u"V;u"V;u"V;u"V;u"V;u"V;u"�
t�+� ��v;/-38X>7vgh4^+X�h�.� JF�0;9fL�0;3fZ�he��V��t.�	�xfnt.XsJv.;u"6����h�_8_�	f�t�;u"'�	�xfnt.XsJv.;u""f�<�tfy�y�t<Xw<	�x.nt.fsXvf;u"&�	�xfnt.fsJv.;u"�(�6�f�r�ٟp��tg�r�ٟ�t`�s�	�xfnt.XsJvf�uh�&�r ?�r��u�r�u�$;u =�t�rXt��u$�r�u��$�J�0��&&�s���pvf;u"��i:�GM�s ��tu�s����s<��t�K;getY�s����9�sf�t,�+M�s���pvf;u =�t�sft���s�;u"V;u"V;u"����hHK�v���nֿ���r.����r.�t��r.���t�rX�u�$�u�$�F�r��u�,�u���\�i;�rft�	�x.nt.Xs<vf;u"���t�,N��~�[���~.�t�~X?��t�M91G�~�;uhV�';u"�z$�2. Jf M U ? > L d
u-/3�;Y���8��[N<2.�n M-�H>�� � i�n���;Kn����|t|>:Me����$<�S��W/j:>�� �}<�<�}t�<�~<K��������u-Ki	� ;�=W=�~t�� �hu����}fLX#.X��LV=;/eL�?�_�J����=-=$�g�g�n.�ge�<Lg��Ek>K� ��� �/�=W=G � �a m 2���~����Z(���}%=s=��l	t� =-=u��L�u� ���x2#��u;K�t.����=-=���~8� �l��g��������u-Ki	� ;�	t��q<��������u-Ki	� ;�	t��q<��������u-Ki	� ;�	tE'�~.�X�~�g��������u-Ki	� ;�	tE8�=-�~��hu-/h�r#�hu-/h�r)�h�ؑr��h�ؑ���=-=�~�g�=-�n<�ge�<�~.�Jh���Ȓg$�g�=-�n<�ge�<�~.�Jh����g�=-�n<�ge�<�g��Ȓgnt��gtu��v�i.�~Ȣg�=-�n<�ge�.�g����=-=� 0aX.? C��ב闑�z�4LV�=-g��T./�K���� X/�=-=��� XaX.? "<e.��ב�t.���z�@�T�/�KfLV�=-g��~֒��/>(���~1V%�u���taX.? C��ב闑�z�4LV�=-g���.hX���/>(���~%g���L� ���xS�LV=;/eL�?$���ב闑�z�~C���/>(���%uZ�� ���x�~'#�u�/�=-=%&a���~f�����0����~;g���Lz�g���L� t��xv#� ��=W=x�g�~t#X��u�i=W=x�g�~t�Xt�#���~�#X��u�i=W=x�g�t� ���=W=x�g@t=W=H�� #�~.�XH�� �w��~.�Xt�~�� ��/ʈx+���I�`�<�.��n�w��~.�X�t�7�=W=��=W=H�7=W=��=-=u��L7t� ��~#� ���� B�~X�pK��<>�~t=��������u-Ki	� ;�	tE�#nhu����}<KW/j:v�El#���=-=$�g�u�nX�ge�<Lg��� 0�}<. �P��.�}<2�� �LV�=-g�?(C���u;/����z�~O/�=-=s2f,=-� ��^(�.���/>�>x@���~/=-=uu;/�L� t��xJ%� .?���tl�� ��~��X�~t��=s=��=W=>�=-��=-=��F��}J�=^��:0�r��<>�|t�<K��������/�=s= �}& ? + ? ����>�u-=i	� ;�Ȅ�������u-/i	� ;�	tE,�3�֦hu-/h���~.�g�=-�n<�ge�<Lg��at�?�_��ב�Yh��~@u�<�~��� �>V=;/eL��~���g��������u-/i	� ;�	tEJZ(���|9��20���g���L� t%��g� $=-=�o��`�l�g�hu-/h�� )�~.g��������u-/i	� ;�	tE�~.g��������u-/i	� ;�	tE�~.g��������u-Ki	� ;�	tE�~��X�~�u���=-=-�g�=-�n<�g�f�g���hu-Kh�� '�~�Ȓg�.=-�~��g�g�n.�g�f�~.�Jhg���#�hu-/h�r#�hu-/h�r)�hu-/h�k#u��ht�=W=�~��#�u���~�Y=sg
�
<?$����t.���z�~BȒgn$Ȓgn$Ȓg$�g�g�n.�g�f�g��a .�~�Z��/�4���~/�g�g�n.�g�f�g���g�g�n.�g�f�g��/�K^(u���~t�� �Y�
t
<?${���闑�z�B���u���~tu���~t/K�KA*=-=u��L� ta .�~�Z���v,���~1� ���x�~�� ֑�
�
t?$����t.���z�D���g���L� �a .�~����/�4���~1� �Y�
t
<?${���闑�z�@��a�.�~�Z���v,��L/���� �/�K(/�K(/�K%.a .? ���闑�z�B����xS�Y=sg
�
<�~�Z��/�4��u/�~.g���L�t.���~��X�����g���L� t��� '��xs���x��g���L� �咈x�~��Xt��n�[�!X�~)�Xt[�!��~)���~.�X�^�=W=\�� �=W=x�g�tO�� '=W=�5������ �=W=x�gw�=W=x�g@t=W=��� �=W=�#	.��� ��#4���~.�Xt��n�����#X�t�~J�X1=W=x�g@t=W=1������ �%)�~f�tgz=W=�~�t�y4�u#��X>�~tK��������u-/i	� ;�	tE�z.�<�y<" t �� X2�}��-/0k)6uMW
X�	JL�g�vf�J�}��I==g�=-=��	���g�x����|tK�XiK�݅��-/
X��}�=-=��~���X=-=��g � g��?+?Y-/fu��}JL�=-=��=-=��=-=�U�K���9M�ht� %=-=���s��f�t�hge�<�
��u<g�
<h=�u;K!��	���g�v<�	.�v<�t��ge�<�g�tK�sX�ge�<�g�tK�sX�ge�<�g�tK�sX�ge�<�g�tK!X�r��ge�<�g�tK^X��s��ge�<�g�tK�rX�ge�<�g�tKtX�sX�ge�<Kg�Y�"Y � � �	 ��t.?+?T��}t)O f��>�~tK��������u-/i	� ;�	tE�|.�.�|<g��:==K�utu�
�G====�v����hu-/h���~���=-=,�g�=-�n<�g�f�;�֦hu�!�z%�	J��g�|����=-="u���|<�t֢g�=-�n<�g�f�g��a .? {���闑�z�~@/�K(Y�
t
<�~�Z���v,��L/���u���~t#Y�
t
<?�{���闑�z�~@=-=u��L� t��x@�/�K�(�� �a .�~�Z���v,��L/����x+�������]��X��~.=-=u��L7t�� �w�3%#�=W=x�g�~t�X�!֡=W=x�g@t=W=1���I�L�7�=W=�!��~#�|-
tz<�K	*/W/u.<s<Kv�iuJ.sJ�u��g
�{=Xy.	JuMLm�lu-/����. of # 9 ? >j����s<.  i�x�tN � � I = = W K��xt�gH<8.;I<���xXV�f�W*'�gMvfM+�Zdh t �i=�yf�.V�wAV>�v;=.�xJ��e�<�g�<�} �g���
���X?+>�u�k��ge�<M+<Tf,tY��p�)�w�}�=-=Yz lz.��u-/ .�.?+>�-Yi�+?Y�k��ge�<�=� <�f� thg�t ���"��{$hu-/0��<�{.Z�=�g-g��-�<<it�uX�
f�ufhgel<B=Hv�
<ytq{W���vX�	f�vf0geYJ�=Hv�
�qqq�w��t�yJ�?��?+?v:0�p�f.D�<��f� �?�?u-/3!J_.*JR
��;�gg�����T�XtvY�u;/����g�ofO�h�s<.��V$g.8Ny<5����g�o�t�"�Ȅ�g�o.�,0%XO73`Jy��s��g�	���i�	Ju-//��pf��=-=Y-/ju-//�k��ge�<Lg=�X�p.�t�p��t=-=��p�-=i�KI@�G�<��h&�,0!�g�<�s<� �728X\ATk;T^<W<).���� ��~X�{.�<<��Jh�y*� .�� h�z*x<��.Y��s<=�J�;M�>,2*@j�=L�9J� �0�'0��$>'$y"q"�Y��,>[K]�>
$#$�"=-=�=-=�/"N"�"�x��ge�<M3<>J<4f����~$��	Jwg����tu����~����u-/i	�   ;�	tE ��jg�u�n��ge�<�g � ��=-=� $>Vg=-g��~�Z��/> �>���0/�=s=�)91 �~���X�~t���~t� �a .?�C���u;/����z�~KN0=-=uu;/�Lt=-� ���=W= y���xV%l�� 䑑e��~��X�~t���=-_�%#�=-= ��F��f�fq<f�	<w.K-E�<.fD<h�n7<D<l�7f/;uN<��.�T<�+�V.4�vt/	.y<gl�ZJ�%J�Z���%'�zf4X�q�flXugutsf=buyvp<y<uvuuvZhr� <��t� <.u.>	<uX.x.D�XY;�� ���@��y.�z.�z�KW�[��$X82[X�[�hd>Vhxp2�K;���I=�;�P/-�Y�m �f�m.�.I=�;�l<e=-g�&tt�Q��g0.���otu����Z�K;9�J�>�
�Ki;/^�L[h.w�rf����� �{�j9�<����x�     �   �      ../../../gcc-4.9.1/libgcc /opt/MeetiXOSProject/MXlibraries/include/eva  libgcc2.c   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   libgcc2.h     ��
�}f�J�}�s.u.0�g����~tX= �ZH0�-0;-L-LIK��L,>)��=� .�~��J�}��f�t -   �   �      ../../../gcc-4.9.1/libgcc /opt/MeetiXOSProject/MXlibraries/include/eva  libgcc2.c   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   libgcc2.h     P��	f�}XKRKMt..0Nf�J�~�J=
Xt� ��~<g��� t�J��Z,0,h�I0,KK-KK-/�+/-/LH0/L)ML��/-��� f�� G   �  �      ../../../gcc-4.9.1/libgcc /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva ../../../gcc-4.9.1/libgcc/../gcc/config/i386 ../../../gcc-4.9.1/libgcc/../include . /opt/MeetiXOSProject/MXlibraries/include  unwind-pe.h   unwind-dw2.c   unwind-dw2-fde.h   unwind.inc   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   i386.h   dwarf2.def   unwind.h   unwind-dw2.h   string.h   stdlib.h     ���]* � u u ; 1M XY�>�.\<q.@��zf�<�z������~<�t�~���t�l�73 xfY�z������~��y.@�.�y<�.�y��uu;1���>u�>:>/i��y ��~X�y uu;1�fg�~X�y�w�,�~�	���u;�Zu;�Z=;0iX�y uu;1y�*5uu;1��ʼu_t�y�uu;1�J�U��y�uu;1�J�G��y�uu;1�J�N��y�uu;1uf2*5uu;1���u|˕���� <\=�gK?9�f� <�X�y�uu;1�f�xX*�.�xf�uu;1�f���X�y�uu;1�f���X�y�uu;1�f�[�xf*�.g�x��uu;1��/�~X�y�uu;1�f�u�x.@*�uu;1���~t�y�uu;1���ʼu�~t�yXuu;1�fY;gZ=��g[�0�~X�y�uu;1y�*5uu;1��ʼu�~t�y�uu;1���ʼu�~t�yXuu;1�f�u�w.@*�uu;1���~t�y�uu;1u�21uu;1�f��Wu�xt=<iu-I0����zX=�~X� �KgX��uu;1� ���KT������J�f3S373EA��uv�w��X�w����V0f�y<�<�wf��u/�yJQ
f���w�uu;1�fIi,uK-g�}tuu;1�JmE]t(��~��Q
J�cȅL�f5X�y�!�	��|<�.�|J1�.�~��X�}t	f������� J���w<�f�wX�J\�vt��	"L�wJuu;1�Jr0�v��7�~�	��'�~��.;=H X�}�uu;1�JvrMf�J��x<=<i�0�<�~�=�~X� KgX� uu;1� ��ItK�/;.i�0��I/@[�w<�f�wX�Jv�w�/;SJ�Xuu;1� J=;zt��=;��yt5x��v��� <h��h�:�0�}�����}th��h��}���my.�M�.�~J���~�k73� %H=��Y �|��f��z��<I=*f�|<\q�vH>����|�� �LI=zXLI=zXLI=zXLI=�X�\:�('�}J�./�~��|J��6���}<�X�}J	f�+�|�uu;1� J�rs�H>���f����|<�s�H>���.��=sKK�~J�.p�IuWK�d1������z<�J=FN����A:L9M�"�==rLK���~J�.�~�=XJ(.�t�K�~.�.���� J�~�|�uu;1���|�uu;1�J�|��s�H>���.��K�~.�.s���~t�.�}X�~.=<��0��t�{�uu;1�fK�{X=���~��|t�� �>H=/���~.�f�.]�{��f.X�}J�./7X�}<�.Z�}.�.Z�}.�.Z�}.�.Z�}.�.Z�}.�.Z�}.�.`�}��.XX�}.�.Z�}t�.Z�}.�.Z�}f�./&X�}��.sX�}��.`�}��.sX�}��.`�}��.�zX��Kr�Kg��<uu;1���q2Zzt5�./W/-I��wf��K��	��uJ*�
.�v�uu;1�
f|��a�]�$t\t<f,��wf�u �t�v��Ii�
t\t�u.*�uu;1�
f�v.�u�	�
X�u.*�uu;1�
f�v.Lu�t�w�wJ	J���wfgu����Lj��	<�v���L�	���v�]t�
t�v����wJ/��	t4zX4z<Pz.lkHwt�x*@u
J�~� ��n��vp�J�wJ/K�	J*���v��	<y��f!`�v�\G�>2xX�
t>zfz�v��~��v��Lg����<�t<�<�s.�JlfXWY zX� �ɭtv����
X�u����v�/`  Xs���u< �
��UKIK>/$�}����}t�t�}<�w.�J�wJ/K�
�u i()��u.�
�tc
��u@�
f�t�Gu>���.km��t.�
�\G�>2 xX �tz�4�u��[H�6:> u. �vtz l5�u�K�~J�f/=��u�u��!u M;�u�u��3)%Sk)y1vq�,v�l	Jt��K-K4wt����u�e/a�.���t�ya&eSk�#Pv��]i��Z!Xd�Xw��<�sfe�� t���sJi;uY[(e==&xb$=e*j�dy�=��\��e=#xb$=a�8�=eu\ XV��e=%���e�Zd0� Xy�
��e=�<Ku�{\�j�\s��;/fq<X�Y `   �  �      ../../../gcc-4.9.1/libgcc /opt/MeetiXOSProject/temp/build-gcc/gcc/include /opt/MeetiXOSProject/MXlibraries/include/eva ../../../gcc-4.9.1/libgcc/../gcc/config/i386 . /opt/MeetiXOSProject/MXlibraries/include  unwind-pe.h   unwind-dw2-fde.c   unwind-dw2-fde.h   stddef.h   stdint.h   kernel.h   fs.h   ipc.h   kernquery.h   i386.h   unwind.h   gthr-default.h   string.h   malloc.h   stdlib.h     ��]* � u u ; 1M XY�>�.�h��.f�2[�ytH	Jw<
.z. �H�fNFR8
< u W = Ո " u ; u ���|X�M	<wX.t Jw<	XI�y<_r�.���M
�@r��t��w<	.z�B��<q.J	f)�g<LY�0g2hm.g=vtu=kf�I1k���uu;1� �u=fH�� t�J=/� <0� �fM=;/Y�#��4z<�IKng  .�~�@�f�I/�~f@�f�~t@�fRxJ�Op<<t<MO�x<x�<Y�=W f�	����gJ�m��|��X�uWKh=Z�M{�iU/�|J�.MYY�|<4�f.�Ke�0b<XMJ7<�H�-uv,"J`J �`JX�}�K�}��f�w�{f�Xi�-/�JݭiU/�{��f3.� �Z,<>�v,%J]J#�]JX==,KK.�z��f�w�z��Xiu;/�J�;�^uiU/�%82�/�|�f�~��fO<0X�~��fK<4Xل#��?GM��� 0gM?Hvyf=I/M?Hvyf,� J.�}fg-Kh�=y)�uXWuK������� ����)�w9�ot؃I/�yJ�f�X�{t�.i9Z:M��~��;Kf/�}t�K;ui;u�t��;=��~�Ke3h�~�	tw.	J6u�2�Oog�">��=K,h�9M0�r<�IA7/N�"�|��$r�gI1)u� t=�Y�u��YK,K���LH',L/t��>�}����#dt�~t� t5�}��~t�J�~��|t�L JjL>Wpg=MRgtf<@�h.�>WuRsfgute��Nic�WpkRgs<uu<e<	.LH�=LuEh=McDge=mpJJq�uKcDufgu
te=f�itKuKzfgvDwf
te<��O � �� e |�� q�f[	X_���Z<&.m�=;/�t`f$���Lyf���.
 vf
J <�L�-/ .�h�I=�y.�f�X=;��b��+=0r.�=-gw� I�+=0 getenv FS_READ_DIRECTORY_EOD FS_TASKED_DELEGATE_REQUEST_TYPE_READ FS_NODE_TYPE_ROOT FsClonefdStatus FS_LENGTH_ERROR FsCreateNodeStatus FS_SEEK_CUR MESSAGE_RECEIVE_MODE_BLOCKING FS_TELL_SUCCESSFUL GET_WORKING_DIRECTORY_ERROR FS_TRANSACTION_NO_REPEAT_ID FS_TASKED_DELEGATE_REQUEST_TYPE_READ_DIRECTORY GET_WORKING_DIRECTORY_SUCCESSFUL MESSAGE_SEND_STATUS_EXCEEDS_MAXIMUM FS_LENGTH_SUCCESSFUL mblen FS_READ_ERROR FS_PIPE_ERROR FS_CREATE_NODE_STATUS_FAILED_NO_PARENT ThreadPriority FS_DIRECTORY_REFRESH_ERROR FS_TRANSACTION_FINISHED wchar_t MESSAGE_RECEIVE_STATUS_EXCEEDS_BUFFER_SIZE FS_NODE_TYPE_MOUNTPOINT FS_CLOSE_SUCCESSFUL MessageReceiveMode SET_WORKING_DIRECTORY_ERROR MESSAGE_SEND_MODE_NON_BLOCKING FS_READ_BUSY FS_WRITE_BUSY FS_TRANSACTION_REPEAT KernqueryStatus FsTransactionID FS_OPEN_NOT_FOUND FS_DISCOVERY_ERROR mbtowc FS_LENGTH_NOT_FOUND MESSAGE_SEND_STATUS_QUEUE_FULL FS_WRITE_SUCCESSFUL FS_SEEK_SUCCESSFUL long long unsigned int FS_DIRECTORY_REFRESH_BUSY FsOpenStatus FS_OPEN_BUSY FsRegisterAsDelegateStatus FS_TRANSACTION_WAITING FS_CLONEFD_INVALID_SOURCE_FD FsSeekMode FS_WRITE_ERROR FS_DISCOVERY_SUCCESSFUL FsNodeType /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/libsupc++ FS_CLONEFD_ERROR THREAD_PRIORITY_NORMAL bsearch FS_READ_INVALID_FD FS_DIRECTORY_REFRESH_SUCCESSFUL free MESSAGE_RECEIVE_STATUS_FAILED_NOT_PERMITTED FS_SEEK_END FS_TELL_INVALID_FD FsDiscoveryStatus FsLengthStatus FS_CLOSE_BUSY FS_LENGTH_INVALID_FD MESSAGE_SEND_MODE_BLOCKING FS_OPEN_SUCCESSFUL SET_WORKING_DIRECTORY_NOT_FOUND ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/del_op.cc 5div_t THREAD_TYPE_VM86 MESSAGE_RECEIVE_STATUS_QUEUE_EMPTY FS_NODE_TYPE_FOLDER FsSeekStatus FS_CREATE_NODE_STATUS_CREATED FsWriteStatus KERNQUERY_STATUS_SUCCESSFUL uint8_t quot FS_LENGTH_BUSY FS_READ_SUCCESSFUL mbstowcs FS_OPEN_DIRECTORY_SUCCESSFUL long long int _ZdlPv FS_NODE_TYPE_FILE FS_CLOSE_INVALID_FD THREAD_PRIORITY_IDLE ThreadType FS_TASKED_DELEGATE_REQUEST_TYPE_DISCOVER THREAD_TYPE_SUB FsPipeStatus ldiv FS_NODE_TYPE_PIPE srand FsOpenDirectoryStatus FsTransactionStatus FS_OPEN_ERROR FS_TASKED_DELEGATE_REQUEST_TYPE_GET_LENGTH THREAD_TYPE_MAIN FS_SEEK_SET MESSAGE_RECEIVE_STATUS_SUCCESSFUL operator delete SET_WORKING_DIRECTORY_NOT_A_FOLDER FS_OPEN_DIRECTORY_ERROR FS_NODE_TYPE_NONE GetWorkingDirectoryStatus FS_CLONEFD_SUCCESSFUL FS_WRITE_INVALID_FD FS_SEEK_ERROR FS_WRITE_NOT_SUPPORTED FS_SEEK_INVALID_FD MessageSendMode MESSAGE_SEND_STATUS_SUCCESSFUL FS_PIPE_SUCCESSFUL FS_CREATE_NODE_STATUS_UPDATED short int FS_TASKED_DELEGATE_REQUEST_TYPE_CLOSE MESSAGE_RECEIVE_STATUS_FAILED FS_REGISTER_AS_DELEGATE_SUCCESSFUL GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=del_op.lo FS_OPEN_DIRECTORY_NOT_FOUND FS_REGISTER_AS_DELEGATE_FAILED_DELEGATE_CREATION uint64_t FsTellStatus FS_READ_DIRECTORY_SUCCESSFUL FS_CLOSE_ERROR FS_READ_DIRECTORY_ERROR MESSAGE_SEND_STATUS_FAILED MESSAGE_RECEIVE_STATUS_INTERRUPTED sizetype strtoul MessageSendStatus KERNQUERY_STATUS_UNKNOWN_ID unsigned char FS_TASKED_DELEGATE_REQUEST_TYPE_WRITE strtod strtol FsReadDirectoryStatus FsReadStatus 6ldiv_t FsCloseStatus FsDirectoryRefreshStatus short unsigned int GET_WORKING_DIRECTORY_SIZE_EXCEEDED atof atoi atol FS_TASKED_DELEGATE_REQUEST_TYPE_OPEN FS_REGISTER_AS_DELEGATE_FAILED_EXISTING FsTaskedDelegateRequestType SET_WORKING_DIRECTORY_SUCCESSFUL system SetWorkingDirectoryStatus FS_DISCOVERY_NOT_FOUND FS_DISCOVERY_BUSY MESSAGE_RECEIVE_MODE_NON_BLOCKING MessageReceiveStatus qsort __unexpected languageSpecificData terminateHandler _ZN10__cxxabiv112__unexpectedEPFvvE _Unwind_Sword unexpectedHandler __cxa_dependent_exception __is_dependent_exception handlerSwitchValue new_ptr check_exception_spec __get_exception_header_from_obj lpstart_encoding cs_lp __is_gxx_exception_class _sleb128_t _Unwind_Context actionRecord __cxxabiv1 __in_chrg TType _URC_FATAL_PHASE1_ERROR _URC_HANDLER_FOUND _Unwind_Exception handlerCount __gxx_dependent_exception_class _URC_NO_REASON ar_disp __get_dependent_exception_from_ue nextException catchTemp get_ttype_entry xh_lsda do_something found_something _Unwind_GetRegionStart _ZN10__cxxabiv111__terminateEPFvvE _URC_END_OF_STACK exc_obj action_table landing_pad __get_object_from_ambiguous_exception _Unwind_Action read_sleb128 saw_cleanup ip_before_insn thrown_ptr _Unwind_Exception_Class filter_value unaligned new_xh _ZSt9terminatev __builtin_unwind_resume private_1 private_2 read_uleb128 adjustedPtr uncaughtExceptions GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=eh_personality.lo _Unwind_Ptr unwindHeader __cxa_exception language_specific_data this p_or_d exceptionDestructor 19_Unwind_Reason_Code action_record __cxa_allocate_exception __get_object_from_ue lsda_header_info _Unwind_Exception_Cleanup_Fn cs_action _Unwind_GetIPInfo _Unwind_SetGR _uleb128_t restore_caught_exception size_of_encoded_value ttype_base ar_filter cs_start _Unwind_GetDataRelBase __terminate catch_type ~end_catch_protect _Unwind_SetIP __cxa_end_catch _URC_NORMAL_STOP ttype_encoding _URC_INSTALL_CONTEXT _ZSt10unexpectedv exc_obj_in LPStart _throw_typet __gxx_primary_exception_class handler_switch_value found_handler __cxa_begin_catch ue_header actions ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/eh_personality.cc exceptionType __cxa_call_unexpected cs_len empty_exception_spec install_context end_catch_protect_obj parse_lsda_header base_of_encoded_value _Unwind_GetLanguageSpecificData __cxa_call_terminate __padding _URC_CONTINUE_UNWIND thrown_ptr_p __cxa_get_globals_fast found_type call_site_encoding primaryException _Unwind_GetTextRelBase get_adjusted_ptr bad_exc _Unwind_Resume _Unwind_Internal_Ptr found_terminate __cxa_eh_globals throw_type _URC_FOREIGN_EXCEPTION_CAUGHT found_cleanup found_handler_type xh_switch_value read_encoded_value_with_base found_nothing xh_terminate_handler __gxx_personality_v0 _URC_FATAL_PHASE2_ERROR saw_handler read_encoded_value save_caught_exception __cxa_throw __cxa_rethrow __get_exception_header_from_ue operator new [] _Znam operator new ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/new_opv.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=new_opv.lo _Znwm decltype(nullptr) ~exception_ptr dest __max_align_ld __max_align_ll GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=eh_throw.lo __gxx_exception_cleanup _ZSt13get_terminatev __get_refcounted_exception_header_from_obj _M_exception_object 11max_align_t referenceCount _ZNSt15__exception_ptr13exception_ptr4swapERS0_ tinfo __cxa_refcounted_exception __exception_ptr _ZNSt15__exception_ptr13exception_ptraSERKS0_ __cxa_get_globals __get_refcounted_exception_header_from_ue operator= _M_addref _ZNSt15__exception_ptr13exception_ptr10_M_releaseEv _ZNKSt15__exception_ptr13exception_ptr6_M_getEv _ZNKSt15__exception_ptr13exception_ptr20__cxa_exception_typeEv nullptr_t _Atomic_word _Unwind_Resume_or_Rethrow operator bool __cxa_exception_type _Unwind_RaiseException _M_get _ZSt14get_unexpectedv get_unexpected ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/eh_throw.cc _ZNSt15__exception_ptr13exception_ptr9_M_addrefEv _ZNSt15__exception_ptr13exception_ptraSEOS0_ _M_release _ZNKSt15__exception_ptr13exception_ptrcvbEv get_terminate __cxa_free_exception GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=eh_call.lo ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/eh_call.cc lconv _S_showpoint _ZNKSt8numpunctIcE8truenameEv __io _ZNSs12_M_leak_hardEv not_eof _S_ios_iostate_end _ZNSt6locale5_Impl16_M_add_referenceEv iostate _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKa _ZNSolsEPSt15basic_streambufIcSt11char_traitsIcEE _vptr.basic_ostream _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKh _ZNSt8ios_base4setfESt13_Ios_Fmtflags _M_install_cache _ZNKSs8capacityEv _ZNSo6sentryD2Ev _ZNSs6resizeEmc __ops _ZNKSt15basic_streambufIcSt11char_traitsIcEE5epptrEv _ZNSs5clearEv _ZNSoC1EPSt15basic_streambufIcSt11char_traitsIcEE __gnu_cxx _ZN9__gnu_cxx13new_allocatorIcE10deallocateEPcm _ZNKSs4findEcm _ZSt5flushIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ _ZNSs4_Rep7_M_grabERKSaIcES2_ _M_refcopy _Reference _S_ate operator==<mbstate_t> _ZNSs13_S_copy_charsEPcS_S_ _ZNSt11char_traitsIcE4findEPKcmRS1_ _M_refcount _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecb _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecd __ios_type __vtt_parm ostreambuf_iterator const_pointer _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecl _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecm _ZNSo9_M_insertIlEERSoT_ _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecx _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecy _M_check_length pos_type _Category _ZNSo9_M_insertIPKvEERSoT_ __np _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_a _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_c _ZNKSs8_M_limitEmm _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_h __cerb _StateT _ZNSs6rbeginEv _S_id_time _M_impl _S_dec _ZNKSt9basic_iosIcSt11char_traitsIcEE5widenEc _ZNSo9_M_insertImEERSoT_ _M_p __os __pos __out __debug __pf setlocale _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_RKSs _ZNKSs7_M_dataEv fpos _ZNSoC1Ev __fmtfl replace _S_showbase _ZNKSs6_M_repEv _Rep_base __state _S_oct _ZNSsaSEc _M_names _ZNKSs4findERKSsm _ZNSt9basic_iosIcSt11char_traitsIcEE5clearESt12_Ios_Iostate __refs _ZNKSs7_M_iendEv _ZNSs5eraseEN9__gnu_cxx17__normal_iteratorIPcSsEES2_ __ret _ZNSs14_M_replace_auxEmmmc _M_check_same_name off_type _ZNSs5beginEv reverse_iterator<__gnu_cxx::__normal_iterator<char const*, std::basic_string<char, std::char_traits<char>, std::allocator<char> > > > __len pubsync _Setfill<char> _S_internal __streambuf_type _S_empty_rep ends<char, std::char_traits<char> > _ZNSt11char_traitsIcE4copyEPcPKcm _ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEEc _S_eofbit __sb num_put<char, std::ostreambuf_iterator<char, std::char_traits<char> > > __sp int_frac_digits _M_destroy _ZN9__gnu_cxx13new_allocatorIcE7destroyEPc rfind _ZNKSt6locale2id5_M_idEv _ZNKSs15_M_check_lengthEmmPKc _ZNSt8ios_base4setfESt13_Ios_FmtflagsS0_ _ZNKSs6substrEmm _S_construct_aux_2 __rhs _ZNKSs9_M_ibeginEv _S_scientific _ZNSo6sentryC2ERSo _ZNSt6locale5_Impl19_M_remove_referenceEv _ZNKSs4copyEPcmm _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St8_SetfillIS3_E _ZNKSt5ctypeIcE5widenEc operator& operator* operator+ __gnu_debug __put _ZNSs12_S_empty_repEv __ineof _ZNSs6assignERKSs _ZNKSt6localeneERKS_ _ZNSs4_Rep8_M_cloneERKSaIcEm currency_symbol __err _ZNSt6localeaSERKS_ _ZNSs6appendEPKc _ZNSo9_M_insertIxEERSoT_ operator| operator~ to_char_type _ZNSoC2Ev output_iterator_tag __exchange_and_add_dispatch substr _ZNSs6insertEmRKSs _ZNKSs4_Rep12_M_is_sharedEv _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKc __ws ctype<char> _M_refdata operator<< <char, std::char_traits<char> > _ZNSt6locale5_Impl16_M_install_cacheEPKNS_5facetEm _ZNSt15basic_streambufIcSt11char_traitsIcEE10pubseekposESt4fposI9mbstate_tESt13_Ios_Openmode _M_coalesce _ZNSo9_M_insertIyEERSoT_ _ZNKSs13find_first_ofEPKcm _ZNKSs7compareEmmPKcm _M_set_length_and_sharable __fmt _ZNSs4_Rep26_M_set_length_and_sharableEm _ZNSt11char_traitsIcE2eqERKcS2_ _ZNSs9_M_assignEPcmc _S_fixed _ZNSs18_S_construct_aux_2EmcRKSaIcE _ZNSs4_Rep10_M_refcopyEv _S_cur __left _ZNSolsEPFRSt8ios_baseS0_E epptr _ZNSs7_M_copyEPcPKcm _ZNSs13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIS_SsEES2_ _ZNKSs7compareEPKc _ZNKSs16find_last_not_ofEcm _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_S1_S1_ ~sentry _Distance _ZNSolsEb _ZNSolsEd _ZNSolsEe _ZNSolsEf _ZNSt6locale5_Impl18_M_check_same_nameEv _ZNKSs2atEm _ZNSolsEl _ZNSolsEm _ZNSolsEs _ZNSolsEt _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_NS0_IPKcSsEES5_ _ZNSolsEx _ZNSolsEy _M_iend _ZNSspLERKSs _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKc _S_create _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St12_Setiosflags _M_insert<bool> _M_off _ZNSt11char_traitsIcE7not_eofERKi _M_caches uncaught_exception _ZNKSt9basic_iosIcSt11char_traitsIcEE10exceptionsEv ~basic_string _ZNKSt19ostreambuf_iteratorIcSt11char_traitsIcEE6failedEv _M_move int_curr_symbol _ZNKSs7compareERKSs _ZNK9__gnu_cxx13new_allocatorIcE7addressERc iterator<std::output_iterator_tag, void, void, void, void> _M_clone _M_replace_safe _ZNSs6appendERKSsmm _M_ibegin clear _ZNSt11char_traitsIcE2ltERKcS2_ _S_end _ZNSs6assignERKSsmm operator!= _ZNSt8ios_base9precisionEl _ZNKSs8_M_checkEmPKc __builtin_strlen _ZNSt6locale5_Impl16_M_replace_facetEPKS0_PKNS_2idE _ZNKSs17find_first_not_ofEPKcm _ZNSs5eraseEN9__gnu_cxx17__normal_iteratorIPcSsEE __check_facet<std::num_put<char> > _M_grab _S_id_collate _M_is_shared _M_widen_init _ZNKSt9basic_iosIcSt11char_traitsIcEE4goodEv __write<char> _S_empty_rep_storage __sbin mon_thousands_sep _ZNKSo6sentrycvbEv _M_assign _ZN9__gnu_cxx13new_allocatorIcE9constructEPcRKc _S_max_size _ZNKSt5ctypeIcE13_M_widen_initEv _ZNSt15basic_streambufIcSt11char_traitsIcEE5pbumpEi _ZNSt9basic_iosIcSt11char_traitsIcEE4initEPSt15basic_streambufIcS1_E find_last_not_of _M_add_reference _S_boolalpha _ZNSt9basic_iosIcSt11char_traitsIcEE8setstateESt12_Ios_Iostate ~locale operator<< <std::char_traits<char> > _ZNKSs12find_last_ofEPKcm _ZNKSs5rfindEcm _ZNKSs13get_allocatorEv _ZNKSs6lengthEv _S_left _ZNSt6locale18_S_initialize_onceEv _M_insert<long int> _M_copy __vtbl_ptr_type _ZNKSs4findEPKcm _S_ios_fmtflags_end _ZNKSs16find_last_not_ofEPKcm _ZNSt11char_traitsIcE11eq_int_typeERKiS2_ _ZNSt15basic_streambufIcSt11char_traitsIcEE7pubsyncEv _ZNSs4_Rep10_M_disposeERKSaIcE _ZNSs6appendEmc _ZNKSs5c_strEv __prec _ZNKSsixEm _ZNSs4_Rep10_M_destroyERKSaIcE _ZNSo9_M_insertIbEERSoT_ _ZSt21__copy_streambufs_eofIcSt11char_traitsIcEElPSt15basic_streambufIT_T0_ES6_Rb _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKcm _ZNKSt8ios_base9_M_getlocEv _ZNSs2atEm _S_badbit _ZNKSs11_M_disjunctEPKc _ZNKSs6rbeginEv reverse_iterator<__gnu_cxx::__normal_iterator<char*, std::basic_string<char, std::char_traits<char>, std::allocator<char> > > > _ZNSt19ostreambuf_iteratorIcSt11char_traitsIcEEppEi _S_out _ZNSt19ostreambuf_iteratorIcSt11char_traitsIcEEppEv _S_right basic_ostream<char, std::char_traits<char> > _M_limit _ZNKSt6localeeqERKS_ pubseekoff _ZNK9__gnu_cxx13new_allocatorIcE8max_sizeEv _ZNSolsEPKv flush<char, std::char_traits<char> > _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKcS4_ _M_replace_category _M_write openmode _ZNSt11char_traitsIcE6lengthEPKc _ZNSt11char_traitsIcE12to_char_typeERKi _ZNSs6appendERKSs _ZNKSs12find_last_ofEcm _ZNSspLEPKc _ZNKSt8numpunctIcE13decimal_pointEv operator[] operator std::streamoff _ZNSt11char_traitsIcE3eofEv _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St8_Setbase _M_insert<long long int> _ZNKSs3endEv _ZNSo9_M_insertIdEERSoT_ __val _ZNKSt4fposI9mbstate_tEcvxEv _ZNKSs4findEPKcmm _ZNSt6locale5_Impl21_M_replace_categoriesEPKS0_i _ZNKSs13find_first_ofEcm __copy_streambufs<char, std::char_traits<char> > allocator_type _ZNSs3endEv __num_put_type _M_insert<double> _ZNSt6locale11_M_coalesceERKS_S1_i _ZNSs6insertEmmc _ZNSs7replaceEmmRKSsmm _ZNSo9_M_insertIeEERSoT_ _ZNSt15basic_streambufIcSt11char_traitsIcEE10pubseekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _M_insert<void const*> _ZNSt6locale5_Impl16_M_install_facetEPKNS_2idEPKNS_5facetE _S_skipws _S_hex _ZNKSs8max_sizeEv _ZNSs6insertEmPKcm _ZNSt11char_traitsIcE6assignERcRKc _M_mutate _M_remove_reference char_traits<char> good _ZNSs6assignEPKcm _ZSt4endsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ _ZNSt4fposI9mbstate_tE5stateES0_ mon_grouping _ZNSs7replaceEmmmc _ZNSs6insertEmRKSsmm _ZSt4endlIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ streamsize find_first_not_of _ZNSs7_M_leakEv _M_leak _M_c _ZNKSs5beginEv _ZN9__gnu_cxx13new_allocatorIcE8allocateEmPKv _ZNSt6locale2idaSERKS0_ _ZNKSs12find_last_ofEPKcmm _ZNKSs5rfindEPKcm _ZNKSt4fposI9mbstate_tEmiERKS1_ ptrdiff_t _Pointer _M_replace_aux __mask _S_floatfield _ZNSt4fposI9mbstate_tEpLEx _ZNKSs5emptyEv append __throw_bad_cast __way _ZNSs6assignEmc _M_insert<long long unsigned int> _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St13_Setprecision _ZNSt9basic_iosIcSt11char_traitsIcEE4fillEc _ZNSs6insertEmPKc _S_id_messages ~basic_ostream _S_facet_categories _ZNSo5writeEPKcl seekp _M_rep _ZNSt19ostreambuf_iteratorIcSt11char_traitsIcEEdeEv _ZSt18uncaught_exceptionv operator&= _S_in _S_initialize_once ~new_allocator _ZNKSs4dataEv _ZNSt11char_traitsIcE4moveEPcPKcm _ZNSs7replaceEmmPKc tellp _M_data _ZNSt11char_traitsIcE6assignEPcmc _ZNSt15basic_streambufIcSt11char_traitsIcEE5sputnEPKcl _ZNKSs17find_first_not_ofEPKcmm _ZNSolsEPFRSoS_E iter_type ~_Alloc_hider eq_int_type _ZNKSt9basic_iosIcSt11char_traitsIcEE7rdstateEv _ZNSs4_Rep9_S_createEmmRKSaIcE _ZNKSs7compareEmmPKc _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_S2_S2_ do_widen _M_base __lhs _ZNSoD1Ev _ZNSs4rendEv _ZNSo5tellpEv to_int_type int_p_sign_posn _S_uppercase GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=ostream-inst.lo _ZNSs4swapERSs _S_classic __normal_iterator<char*, std::basic_string<char, std::char_traits<char>, std::allocator<char> > > __sbout _ZNSs6appendEPKcm mon_decimal_point _ZNSt6locale6globalERKS_ streampos _ZNSo5seekpESt4fposI9mbstate_tE _S_construct __normal_iterator<char const*, std::basic_string<char, std::char_traits<char>, std::allocator<char> > > _M_facets_size _Traits basic_ios<char, std::char_traits<char> > __ostream_type _M_put reserve _ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEEmc rdbuf _ZNSs7replaceEmmRKSs _M_facets __mem __mode _ZNSt11char_traitsIcE7compareEPKcS2_m _S_categories operator+= _M_replace_categories _ZNSoC2EPSt15basic_streambufIcSt11char_traitsIcEE _Alloc operator++ _ZNSs6resizeEm __ostream_fill<char, std::char_traits<char> > ostreambuf_iterator<char, std::char_traits<char> > _ZNSs13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIPKcSsEES4_ _M_dataplus _ZNSsaSEPKc push_back _ZNKSt9basic_iosIcSt11char_traitsIcEE3tieEv _S_terminal _ZNKSt4fposI9mbstate_tEplEx _Rep _M_getloc _M_id pubseekpos _S_ios_openmode_end _ZNSt15basic_streambufIcSt11char_traitsIcEE5sputcEc _ZNSs9_M_mutateEmmm _ZNSspLEc _ZNKSt8numpunctIcE13thousands_sepEv _ZNSolsEPFRSt9basic_iosIcSt11char_traitsIcEES3_E operator-= _M_capacity _ZNSt6locale21_S_normalize_categoryEi _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPKv _ZNSoD2Ev _ZNKSs13find_first_ofEPKcmm int_p_sep_by_space _ZNSs7_M_dataEPc _S_refcount _ZNKSs12find_last_ofERKSsm __ostream_write<char, std::char_traits<char> > _ZNSs12_S_constructEmcRKSaIcE _OutIter endl<char, std::char_traits<char> > const_reverse_iterator basic_string<char, std::char_traits<char>, std::allocator<char> > __dir int_n_sign_posn _S_compare const_reference _ZNKSs5rfindEPKcmm new_allocator<char> _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basece _S_id_monetary _ZNKSs17find_first_not_ofEcm _S_normalize_category _M_length _ZNKSs16find_last_not_ofEPKcmm _S_initialize _ZNKSt8ios_base5widthEv _ZNSt19ostreambuf_iteratorIcSt11char_traitsIcEE6_M_putEPKcl int_n_cs_precedes erase _ZNKSs17find_first_not_ofERKSsm _ZNKSt9basic_iosIcSt11char_traitsIcEE4fillEv ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/ostream-inst.cc _ZSt16__ostream_insertIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_PKS3_l _ZNKSs4rendEv _ZNKSt4fposI9mbstate_tE5stateEv _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St14_Resetiosflags rdstate _M_ok basic_streambuf<char, std::char_traits<char> > _M_set_sharable _M_os ~_Impl __check_facet<std::ctype<char> > _ZNSt8ios_base5widthEl _ZNSo8_M_writeEPKcl _ZNSs9push_backEc _M_insert<long unsigned int> _ZSt16__throw_bad_castv _ZNSt6locale13_S_initializeEv _ZNKSs4_Rep12_M_is_leakedEv seekdir _ZNKSt6locale4nameEv numpunct<char> _S_goodbit _ZNSt4fposI9mbstate_tEmIEx _ZNKSt9basic_iosIcSt11char_traitsIcEE4failEv _S_showpos _S_ios_seekdir_end _ZNSs15_M_replace_safeEmmPKcm _ZNKSs7compareEmmRKSsmm operator- _M_dispose __fill _ZNSs4_Rep13_M_set_leakedEv _S_basefield _ZNSs4_Rep12_S_empty_repEv _ZNKSt15basic_streambufIcSt11char_traitsIcEE4pptrEv _ZNSs13_S_copy_charsEPcPKcS1_ _S_global _ZNSo5flushEv _S_unitbuf _S_trunc _ZNSt11char_traitsIcE11to_int_typeERKc _M_set_leaked fmtflags _ZNSs4_Rep15_M_set_sharableEv _ZNSs7_M_moveEPcPKcm int_n_sep_by_space __off none _ZNSoD0Ev _ZNSsaSERKSs fpos<mbstate_t> _ZNSt9basic_iosIcSt11char_traitsIcEE11_M_setstateESt12_Ios_Iostate _ZNSt6locale7classicEv _S_failbit _ZNSolsEi _ZNSolsEj _ZNKSs13find_first_ofERKSsm _ZNSt6locale5_Impl19_M_replace_categoryEPKS0_PKPKNS_2idE _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St5_Setw _M_replace_facet __c1 __c2 _ZNSs10_S_compareEmm _Facet __wide _ZNKSs4sizeEv _S_id_numeric _ZNK9__gnu_cxx13new_allocatorIcE7addressERKc __ch _S_beg _ZNSs5eraseEmm _ZNSs4_Rep10_M_refdataEv _M_check _S_id_ctype _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_mc const_iterator _M_mask _S_adjustfield _M_install_facet _ZNKSs5rfindERKSsm _M_insert<long double> find_last_of _ZNKSt9basic_iosIcSt11char_traitsIcEE5rdbufEv sputc _ZNKSs16find_last_not_ofERKSsm _CharT _M_sbuf __numpunct_cache<char> localeconv operator<< _ValueT _ZNKSt4fposI9mbstate_tEmiEx __result _ZNSs6assignEPKc _M_state _ZNSs7replaceEmmPKcm _ZNKSt8ios_base5flagsEv _ZNKSt5ctypeIcE8do_widenEc _ZNKSs7compareEmmRKSs __exchange_and_add_single operator== __old _M_disjunct exceptions _ZNKSt8numpunctIcE8groupingEv _M_setstate _S_copy_chars _ZNSs7reserveEm _M_index _ZNSt6locale5_ImplaSERKS0_ _S_bin __copy_streambufs_eof<char, std::char_traits<char> > int_p_cs_precedes _M_failed _M_n _M_is_leaked _M_leak_hard _ZNSt19ostreambuf_iteratorIcSt11char_traitsIcEEaSEc npos ~basic_ios _ZNKSt8numpunctIcE9falsenameEv _ZNSo3putEc /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/src/c++98 __ostream_insert<char, std::char_traits<char> > operator|= _ZNSsixEm ~allocator _S_app _ZNSo5seekpExSt12_Ios_Seekdir find_first_of buffered_bytes_read uint32_t syncungetc _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE8syncputcEi xsputn xsgetn _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED0Ev syncputc _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED2Ev impl_seterr fgetpos ssize_t _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE9underflowEv _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE6xsgetnEPcl _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE9pbackfailEi impl_error impl_reopen _M_file impl_write fclose _M_unget_buf _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE10syncungetcEi syncgetc impl_tell basic_istream<char, std::char_traits<char> > ftell impl_clearerr buffer_size pbackfail file_descriptor fread _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4syncEv ferror ~basic_streambuf _ZSt7getlineIcSt11char_traitsIcESaIcEERSt13basic_istreamIT_T0_ES7_RSbIS4_S5_T1_ES4_ fsetpos buffered_bytes_read_offset ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/misc-inst.cc remove _ZStlsIcSt11char_traitsIcESaIcEERSt13basic_ostreamIT_T0_ES7_RKSbIS4_S5_T1_E underflow _ZSt7getlineIcSt11char_traitsIcESaIcEERSt13basic_istreamIT_T0_ES7_RSbIS4_S5_T1_E setvbuf rename getchar off_t feof impl_eof _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC2EP4FILE __is impl_fileno uflow getline<char, std::char_traits<char>, std::allocator<char> > fopen operator<< <char, std::char_traits<char>, std::allocator<char> > rewind _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE5uflowEv fseek tmpnam buffer_mode stdio_sync_filebuf<char, std::char_traits<char> > _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE8syncgetcEv tmpfile perror GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=misc-inst.lo _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode __str __eof fgetc __c_file fpos_t _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE8overflowEi impl_read impl_close _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE7seekposESt4fposI9mbstate_tESt13_Ios_Openmode buffered_bytes_write __whence fgets _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE6xsputnEPKcl prev impl_seek fflush ~stdio_sync_filebuf freopen _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4fileEv use_facet<std::ctype<char> > __bitmasksize __builtin_memchr operator>><char, std::char_traits<char>, std::allocator<char> > _ZNKSt8ios_base6getlocEv __bit __cdelim snextc _ZNSt15basic_streambufIcSt11char_traitsIcEE12__safe_gbumpEl _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_PS3_ __size __idelim __high ctype_base _ZNSt15basic_streambufIcSt11char_traitsIcEE6snextcEv __low sgetc isgraph __ctype_type _ZNSi6ignoreEli _ZNSt15basic_streambufIcSt11char_traitsIcEE5sgetcEv __safe_gbump ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/istream.cc min<long int> __ct __char_type __bitcur _ZStrsIcSt11char_traitsIcESaIcEERSt13basic_istreamIT_T0_ES7_RSbIS4_S5_T1_E operator>><char, std::char_traits<char> > __large_ignore _ZNSt15basic_streambufIcSt11char_traitsIcEE5gbumpEi _ZNSi7getlineEPclc __testoff _ZNKSt5ctypeIcE2isEjc sbumpc __testis _ZNKSt5ctypeIcE7scan_isEjPKcS2_ _ZNSt15basic_streambufIcSt11char_traitsIcEE6sbumpcEv GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=istream.lo _ZNSi6ignoreEl getline __extracted _ZSt9use_facetISt5ctypeIcEERKT_RKSt6locale isspace memcpy __in __num _ZNKSt15basic_streambufIcSt11char_traitsIcEE5egptrEv __int_type scan_is ispunct _ZNKSt15basic_streambufIcSt11char_traitsIcEE4gptrEv iscntrl __delim _ZNKSi6sentrycvbEv isprint __size_type __s1 __s2 _ExternT __testdecfound operator delete [] _M_extract_int<long int> _Cache _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intImEES3_S3_RSt8ios_basecT_ ~messages_byname _M_find<char> _ZNSt17__timepunct_cacheIcE8_M_cacheERKSt6locale _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecy tm_sec _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm has_facet<std::num_put<char> > _ZSt9has_facetISt11__timepunctIcEEbRKSt6locale _ZNSt7collateIcED2Ev _ZNKSt8messagesIcE8do_closeEi _M_convert_to_char _ZNKSt10moneypunctIcLb0EE14do_curr_symbolEv __sign __k2 __add_unsigned<long unsigned int> _S_destroy_c_locale __dates __adjust _M_extract_int<long long int> __end _ZSt9use_facetISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _M_falsename_size _ZSt17__verify_groupingPKcmRKSs _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNK9__gnu_cxx17__normal_iteratorIPKcSsE4baseEv __tmperr _ZN9__gnu_cxx17__normal_iteratorIPKcSsEmmEi _S_oudigits _ZNKSt11__timepunctIcE20_M_date_time_formatsEPPKc _ZNKSt10moneypunctIcLb1EE11curr_symbolEv has_facet<std::__timepunct<char> > __case_offset _ZN9__gnu_cxx17__normal_iteratorIPKcSsEmmEv _ZSt9use_facetISt8numpunctIcEERKT_RKSt6locale __enable_if<true, long unsigned int> do_transform _ZNK9__gnu_cxx17__normal_iteratorIPcSsEmiEl _ZNKSt8messagesIcE20_M_convert_from_charEPc iterator_traits<char const*> __lc part __lo _ZNSt10__num_base15_S_format_floatERKSt8ios_basePcc do_thousands_sep operator==<char, std::char_traits<char> > _M_day2 _ZSt9has_facetISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _M_day4 _ZSt14__convert_to_vIeEvPKcRT_RSt12_Ios_IostateRKPi time_t __format __newlen __last _ZNSt17moneypunct_bynameIcLb1EED2Ev __mp _ZNSt10moneypunctIcLb0EEC2EPSt18__moneypunct_cacheIcLb0EEm __add_grouping<char> _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _S_iend _ZNSt7collateIcEC2Em _S_get_c_locale _M_time_format has_facet<std::money_put<char> > __basefield _ZN9__gnu_cxx17__normal_iteratorIPcSsEpLEl do_pos_format ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/locale-inst.cc _ZNKSt10moneypunctIcLb0EE11do_groupingEv _ZNKSt8numpunctIcE16do_decimal_pointEv time_put_byname<char, std::ostreambuf_iterator<char, std::char_traits<char> > > _ZSt14__convert_to_vIfEvPKcRT_RSt12_Ios_IostateRKPi _ZNKSt8messagesIcE6do_getEiiiRKSs _ZNSt18__moneypunct_cacheIcLb0EE8_M_cacheERKSt6locale ~numpunct _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcm _ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEEdeEv use_facet<std::collate<char> > _ZNSt18__moneypunct_cacheIcLb0EED2Ev _ZNSt8messagesIcED2Ev __positive_sign no_order __builtin_va_list _M_falsename ~time_put __paddec _M_grouping_size __idx num_get<char, std::istreambuf_iterator<char, std::char_traits<char> > > _M_month01 _M_month03 _M_month05 _M_month06 _M_month07 _M_month08 _M_month09 _M_initialize_moneypunct __conditional_type<true, long unsigned int, long long unsigned int> islower iterator_category _S_atoms_in __plus _M_extract_name __names _ZNSt18__moneypunct_cacheIcLb1EED0Ev __found_zero _ZNSt11__timepunctIcEC2EPSt17__timepunct_cacheIcEm _ZNSt6locale5facet18_S_create_c_localeERPiPKcS1_ _ZNSt15messages_bynameIcEC2EPKcm has_facet<std::time_put<char> > _M_month11 __enable_if<true, int> _ZNSt11__timepunctIcEC2Em _ZNK9__gnu_cxx17__normal_iteratorIPcSsEptEv time_base __builtin_memset _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecl _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _M_extract_num __res _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16do_get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm ~collate_byname _M_c_locale_collate _ZNSt8ios_base5flagsESt13_Ios_Fmtflags _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSs _ZNKSt8messagesIcE7do_openERKSsRKSt6locale _ZN9__gnu_cxx17__normal_iteratorIPKcSsEpLEl _ZNSt7collateIcE2idE _ZSt9use_facetISt7codecvtIcc9mbstate_tEERKT_RKSt6locale __curr_symbol _ZNKSt11__timepunctIcE7_M_daysEPPKc __num_base _S_construct_pattern localtime _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcm _M_day5 use_facet<std::moneypunct<char, false> > _ZSt9has_facetISt10moneypunctIcLb0EEEbRKSt6locale __fbuf __initialize_p __max_digits __width __int_to_char<char, long unsigned int> __sav __builtin_strcmp _ZNSt18__moneypunct_cacheIcLb1EEaSERKS0_ __ctype _ZSt9use_facetISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale __sign_size _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPK2tmcc __only_zeros _ZNKSt10moneypunctIcLb1EE8groupingEv __tm do_grouping __to __tp _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE24_M_extract_wday_or_monthES3_S3_RiPPKcmRSt8ios_baseRSt12_Ios_Iostate _ZNKSt10moneypunctIcLb1EE13thousands_sepEv operator-<char*, std::basic_string<char> > do_negative_sign __first _ZSt9has_facetISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZNKSt10moneypunctIcLb0EE13decimal_pointEv _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe __use_cache<std::__numpunct_cache<char> > _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_bRSt8ios_basecRKSs _M_decimal_point dateorder _ZSt9has_facetISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _S_pad __type time_put<char, std::ostreambuf_iterator<char, std::char_traits<char> > > _M_c_locale_timepunct __ul _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE12_M_group_intEPKcmcRSt8ios_basePcS9_Ri __beg _ZNKSt10moneypunctIcLb1EE16do_thousands_sepEv _M_allocated _ZNKSt10moneypunctIcLb0EE13do_neg_formatEv __found_sci __args collate<char> _M_extract_wday_or_month _ZNKSt10moneypunctIcLb0EE16do_decimal_pointEv __enable_if<true, unsigned int> _ZNK9__gnu_cxx17__normal_iteratorIPcSsEdeEv _M_transform __use_cache<std::__moneypunct_cache<char, false> > _ZNKSt10moneypunctIcLb1EE13negative_signEv __hi2 __date _ZNSt8messagesIcEC2EPiPKcm _ZNKSt10moneypunctIcLb1EE14do_curr_symbolEv use_facet<std::numpunct<char> > __min _ZSt9has_facetISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZNSt14codecvt_bynameIcc9mbstate_tED2Ev _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _M_insert_float<double> __wp _ZNKSt5ctypeIcE5widenEPKcS2_Pc __dnew random_access_iterator_tag _ZNSt15messages_bynameIcED0Ev __matches_lengths use_facet<std::time_put<char> > __declen _M_extract_via_format _ZNKSt10moneypunctIcLb1EE13do_pos_formatEv _ZSt9use_facetISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale __indexlen _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIyEES3_S3_RSt8ios_basecT_ _S_atoms _M_amonth02 _M_amonth03 _M_amonth05 _M_amonth06 _ZNKSt10moneypunctIcLb1EE16do_negative_signEv _M_amonth08 _M_amonth09 _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev clock _ZNSt17moneypunct_bynameIcLb0EEC2EPKcm difference_type _ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPK2tmPKcSB_ _M_insert_float<long double> _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIlEES3_S3_RSt8ios_basecT_ _M_amonth11 _M_amonth12 _ZNKSt7collateIcE12_M_transformEPcPKcm __last_pos _ZNSt17moneypunct_bynameIcLb0EED2Ev _ZNK9__gnu_cxx17__normal_iteratorIPKcSsEmiEl _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev _M_grouping ~moneypunct _M_use_grouping _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _M_curr_symbol _ZNSt15messages_bynameIcED2Ev _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14do_get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _InputIterator __pend _ZSt9has_facetISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZNKSt10moneypunctIcLb1EE13positive_signEv _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_bRSt8ios_basecRKSs __c_locale __days __months2 _ZSt13__int_to_charIcmEiPT_T0_PKS0_St13_Ios_Fmtflagsb __is_null_pointer<char const> __maxlen do_decimal_point __pad<char, std::char_traits<char> > _ZNK9__gnu_cxx17__normal_iteratorIPKcSsEplEl _M_atoms_out catalog _ZSt9use_facetISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Em ~num_put __i2 __i3 _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev __digit __olds _ZNSt8numpunctIcE2idE _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt10moneypunctIcLb0EE11curr_symbolEv _ZNKSt7collateIcE7do_hashEPKcS2_ asctime _S_zero _InternT __convert_to_v<double> __testipad __static_initialization_and_destruction_0 _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev do_narrow isalnum _ZSt9use_facetISt8messagesIcEERKT_RKSt6locale _ZNSt14collate_bynameIcED0Ev has_facet<std::ctype<char> > _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb0EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs _M_extract<true> _ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecPK2tmcc _M_day1 _ZNKSt11__timepunctIcE15_M_time_formatsEPPKc _M_day3 numpunct_byname<char> _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _M_day6 _M_day7 _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv _M_current __days1 __days2 __testvalid messages_byname<char> _ZNSt11__timepunctIcEC2EPiPKcm __add_unsigned<long long int> _M_months __negative_sign has_facet<std::money_get<char> > _M_truename_size _M_date_time_format __member _ZSt24__throw_out_of_range_fmtPKcz _ZNKSt11__timepunctIcE21_M_months_abbreviatedEPPKc _Intl _ZSt14__add_groupingIcEPT_S1_S0_PKcmPKS0_S5_ _M_days __throw_out_of_range_fmt _M_negative_sign_size do_curr_symbol _ZNSt10moneypunctIcLb0EE2idE _M_convert_from_char _M_months_abbreviated _M_date_time_era_format istreambuf_iterator _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _M_date_format _M_days_abbreviated _S_atoms_out _M_atoms_in _ZSt9use_facetISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSs _ZNKSt10moneypunctIcLb0EE14do_frac_digitsEv _ZNKSt8messagesIcE5closeEi _ZNSt8messagesIcE2idE _ZNKSt7collateIcE7compareEPKcS2_S2_S2_ _ZNSt17__timepunct_cacheIcED0Ev _M_group_int _ZNKSt11__timepunctIcE15_M_date_formatsEPPKc __truename operator!=<char, std::char_traits<char> > __ptr _ZNSt17__timepunct_cacheIcEC2Em _Container _ZNSt11__timepunctIcED0Ev use_facet<std::codecvt<char, char, mbstate_t> > do_get_date _ZNKSt10moneypunctIcLb0EE13thousands_sepEv _M_date_era_format _S_clone_c_locale __nskipped _S_create_c_locale _ZNSt16__numpunct_cacheIcEaSERKS0_ _ZNKSt10moneypunctIcLb1EE11frac_digitsEv __matches ~__timepunct_cache _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Em _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm __units _ZNKSt10moneypunctIcLb1EE16do_positive_signEv _ZNSt10moneypunctIcLb1EE24_M_initialize_moneypunctEPiPKc use_facet<std::num_put<char> > _ZNKSt11__timepunctIcE9_M_monthsEPPKc iterator_traits<char*> _ZNKSt10moneypunctIcLb0EE16do_thousands_sepEv _ZNSt17moneypunct_bynameIcLb1EEC2EPKcm __caches _ZSt9has_facetISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale istreambuf_iterator<char, std::char_traits<char> > _ZNSt18__moneypunct_cacheIcLb1EEC2Em _M_time_formats _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNSt6locale5facet15_S_get_c_localeEv _ZNSs16_S_construct_auxIPKcEEPcT_S3_RKSaIcESt12__false_type __xtrc __enable_if<true, long long unsigned int> _ZNKSt8numpunctIcE11do_groupingEv _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE __dat __dt __moneypunct_cache<char, true> __hi1 _M_truename _ZSt14__convert_to_vIdEvPKcRT_RSt12_Ios_IostateRKPi _ZNKSt11__timepunctIcE8_M_am_pmEPPKc _InIter __grouping _ZNSt10moneypunctIcLb0EE4intlE do_open _M_extract<false> _ZNKSt11__use_cacheISt18__moneypunct_cacheIcLb1EEEclERKSt6locale __news _ZNSt10moneypunctIcLb1EE4intlE _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ has_facet<std::num_get<char> > _Cond _M_name_timepunct __found_grouping _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt5ctypeIcE8do_widenEPKcS2_Pc money_put<char, std::ostreambuf_iterator<char, std::char_traits<char> > > _ZN9__gnu_cxx17__normal_iteratorIPcSsEmIEl _M_name_messages _ZNKSt8numpunctIcE11do_truenameEv _M_initialize_timepunct _ZNSt19istreambuf_iteratorIcSt11char_traitsIcEEppEi _M_insert_int<long unsigned int> __sep _S_ominus _ZNSt19istreambuf_iteratorIcSt11char_traitsIcEEppEv __set operator==<char> _ZNKSt10moneypunctIcLb0EE16do_negative_signEv _S_construct_aux<char const*> do_date_order tm_min use_facet<std::money_get<char> > _ZNSt6locale5facet17_S_clone_c_localeERPi _ZNSt16__numpunct_cacheIcED2Ev ~time_get_byname clock_t use_facet<std::time_get<char> > _M_extract_int<long long unsigned int> _ZSt9has_facetISt8numpunctIcEEbRKSt6locale do_get __vend _S_timezones _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_numES3_S3_RiiimRSt8ios_baseRSt12_Ios_Iostate has_facet<std::numpunct<char> > _ZNKSt11__timepunctIcE15_M_am_pm_formatEPKc _ZSt9use_facetISt11__timepunctIcEERKT_RKSt6locale _ZNKSt8messagesIcE4openERKSsRKSt6locale __new _M_positive_sign _ZNKSt10moneypunctIcLb1EE13decimal_pointEv _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb1EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs messages_base moneypunct<char, true> GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=locale-inst.lo isxdigit __cxa_bad_cast _M_am _ZNSt14collate_bynameIcED2Ev __p2 _ZSt9has_facetISt7collateIcEEbRKSt6locale _ZNKSt7collateIcE4hashEPKcS2_ _S_oplus _ZNSs12_S_constructIPKcEEPcT_S3_RKSaIcESt20forward_iterator_tag do_close _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_bRSt8ios_basece _FwdIterator _ZNKSt11__timepunctIcE19_M_days_abbreviatedEPPKc ~collate __moneypunct_cache<char, false> _ZN9__gnu_cxx17__normal_iteratorIPKcSsEmIEl operator() __mult __add_unsigned<short unsigned int> __add_unsigned<long long unsigned int> _ZNSt8numpunctIcEC2EPim _S_iX __valuec _S_ie __unsigned_type money_base tm_wday _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Em time_get<char, std::istreambuf_iterator<char, std::char_traits<char> > > _S_ix __which _ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE9_M_at_eofEv _M_frac_digits _M_month02 _M_month04 __ilen __ps __dfault __wcs __max _ZNSt17moneypunct_bynameIcLb0EE4intlE _ZNKSt10moneypunctIcLb0EE10neg_formatEv _M_am_pm_format __bufend has_facet<std::collate<char> > _M_positive_sign_size __testfail _ZNSs12_S_constructIPKcEEPcT_S3_RKSaIcE do_get_weekday tm_mon __time do_get_monthname _M_negative_sign _ZNSt10moneypunctIcLb1EE2idE _Iftrue _ZNKSt8numpunctIcE12do_falsenameEv _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNSt15numpunct_bynameIcED2Ev __timepunct_cache<char> use_facet<std::__timepunct<char> > _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev codecvt_byname<char, char, mbstate_t> _ZNSt11__timepunctIcED2Ev tm_year _ZNKSt10moneypunctIcLb1EE14do_frac_digitsEv _ZNSt18__moneypunct_cacheIcLb0EEC2Em _M_month10 _ZNSt8messagesIcEC2Em _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _M_month12 _ZNSt15numpunct_bynameIcED0Ev __dynamic_cast ~__numpunct_cache _M_pad __months1 __lit _GLOBAL__sub_I_locale_inst.cc __two _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb0EEES3_S3_RSt8ios_basecRKSs _ZNSt16__numpunct_cacheIcEC2Em _ZSt9use_facetISt7collateIcEERKT_RKSt6locale do_get_year _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev __builtin_vsprintf _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE15_M_insert_floatIeEES3_S3_RSt8ios_baseccT_ _ZNKSt8messagesIcE4openERKSsRKSt6localePKc _ZNSt8numpunctIcE22_M_initialize_numpunctEPi _ZNSt6locale5facet19_S_destroy_c_localeERPi __gbeg _ZNKSt5ctypeIcE6narrowEcc __grouping_tmp _ZNSt18__moneypunct_cacheIcLb1EED2Ev ~time_put_byname _M_amonth01 __distance<char const*> _M_amonth07 __negative _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf _M_aday1 _M_aday2 do_put _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj _M_aday5 _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl _ZdaPv __smax _ZNKSt10moneypunctIcLb0EE13do_pos_formatEv _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy _ZNKSt10moneypunctIcLb0EE13positive_signEv ~messages _ZN9__gnu_cxx17__normal_iteratorIPcSsEppEi _S_oE _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm _ZNKSt7collateIcE10_M_compareEPKcS2_ _ZN9__gnu_cxx17__normal_iteratorIPcSsEppEv _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecPKv _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe __grouping_size _S_oX _M_am_pm _S_oe basic_string<char const*> __cs _Iffalse _S_ox do_frac_digits _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt _ZNSt10moneypunctIcLb0EEC2EPiPKcm _S_iplus _M_insert_int<long long int> _M_amonth10 _ZSt9use_facetISt10moneypunctIcLb0EEERKT_RKSt6locale do_positive_sign _Type _ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE6_M_getEv _ZNKSt10moneypunctIcLb0EE16do_positive_signEv _ZNSt10moneypunctIcLb0EE24_M_initialize_moneypunctEPiPKc operator-> difftime _M_atoms tm_yday _ZNKSt5ctypeIcE9do_narrowEcc __months _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6_M_padEclRSt8ios_basePcPKcRi _M_c_locale_messages _M_extract_int<unsigned int> __lo1 _S_get_c_name _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_bRSt8ios_basece do_compare tm_hour __ws2 do_neg_format __ws3 _S_format_float __name _ZNSt8numpunctIcEC2Em use_facet<std::num_get<char> > __testoverflow _M_compare _ZNSt10money_base20_S_construct_patternEccc __loc has_facet<std::codecvt<char, char, mbstate_t> > _S_iminus has_facet<std::messages<char> > __cloc scan_not _Iter _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE21_M_extract_via_formatES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKc __buf __add_unsigned<long int> __tmpmon _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNKSt10moneypunctIcLb0EE11frac_digitsEv _M_extract_float _S_iE _ZNSt18__moneypunct_cacheIcLb0EEaSERKS0_ tm_mday _ZSt16__convert_from_vRKPiPciPKcz ~numpunct_byname min<long unsigned int> _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Em gmtime _ZSt9use_facetISt10moneypunctIcLb1EEERKT_RKSt6locale __uc _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16_M_extract_floatES3_S3_RSt8ios_baseRSt12_Ios_IostateRSs ~num_get _ZNSt11__timepunctIcE2idE _ZNSt14collate_bynameIcEC2EPKcm _S_minus __cache collate_byname<char> _ZNKSt5ctypeIcE7toupperEc _M_aday3 _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE15_M_extract_nameES3_S3_RiPPKcmRSt8ios_baseRSt12_Ios_Iostate _M_aday4 _M_aday6 _ZNKSt8numpunctIcE16do_thousands_sepEv _ZNKSt10moneypunctIcLb1EE10neg_formatEv _ZNKSt10moneypunctIcLb1EE10pos_formatEv __k1 _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _M_cache _ZNSt10moneypunctIcLb0EEC2Em _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZN9__gnu_cxx17__normal_iteratorIPKcSsEppEi _ZNSt8numpunctIcEC2EPSt16__numpunct_cacheIcEm _S_izero _M_group_float _ZN9__gnu_cxx17__normal_iteratorIPKcSsEppEv operator-- messages<char> _Iterator __qend __dec _ZNK9__gnu_cxx17__normal_iteratorIPcSsEplEl _ZNKSt11__use_cacheISt18__moneypunct_cacheIcLb0EEEclERKSt6locale _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE15_M_insert_floatIdEES3_S3_RSt8ios_baseccT_ __convert_to_v<float> __tm_zone _ZNKSt10moneypunctIcLb1EE11do_groupingEv do_falsename _M_at_eof __value ~moneypunct_byname __found_dec _S_odigits __flags _InIterator isalpha _ZNSt17moneypunct_bynameIcLb1EE4intlE _S_construct<char const*> __gsize _M_pm do_get_time _ZNK9__gnu_cxx17__normal_iteratorIPKcSsEptEv __tmpwday isupper input_iterator_tag _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ use_facet<std::money_put<char> > _S_odigits_end _ZNK9__gnu_cxx17__normal_iteratorIPKcSsEixEl _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev _M_amonth04 _M_extract_int<long unsigned int> _M_insert_int<long int> __mod __oct __priority _ZNSt18__moneypunct_cacheIcLb1EE8_M_cacheERKSt6locale _ZNKSt7collateIcE9transformEPKcS2_ strftime _ZNSt7collateIcED0Ev _M_insert<false> _RandomAccessIterator _ZNKSt10moneypunctIcLb0EE10pos_formatEv __plen _ZNSt7collateIcEC2EPim _M_insert<true> has_facet<std::time_get<char> > _S_oudigits_end __donef tm_isdst _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt10moneypunctIcLb1EEC2EPiPKcm ~__moneypunct_cache __donet _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIxEES3_S3_RSt8ios_basecT_ __lit_zero _ZNKSt5ctypeIcE8scan_notEjPKcS2_ __convert_to_v<long double> _ZNSt14codecvt_bynameIcc9mbstate_tED0Ev _ZSt9has_facetISt8messagesIcEEbRKSt6locale _M_curr_symbol_size _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Em __facets _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE14_M_group_floatEPKcmcS6_PcS7_Ri use_facet<std::messages<char> > __testf _ZNSt15numpunct_bynameIcEC2EPKcm _ZNKSt11__timepunctIcE6_M_putEPcmPKcPK2tm ~money_get _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ iterator<std::input_iterator_tag, char, long long int, char*, char&> _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt __times _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy __uppercase _M_aday7 _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm __fixed __int_to_char<char, long long unsigned int> _ZNSt17moneypunct_bynameIcLb1EED0Ev _ZSt13__int_to_charIcyEiPT_T0_PKS0_St13_Ios_Fmtflagsb _ZNSt6locale5facet13_S_get_c_nameEv moneypunct_byname<char, true> __ampm __verify_grouping __falsename ~__timepunct _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNK9__gnu_cxx17__normal_iteratorIPcSsE4baseEv __msg money_get<char, std::istreambuf_iterator<char, std::char_traits<char> > > _ZNKSt8messagesIcE3getEiiiRKSs __normal_iterator _S_default_pattern do_hash codecvt<char, char, mbstate_t> __oldlen _ZNKSt10moneypunctIcLb1EE13do_neg_formatEv __digits has_facet<std::moneypunct<char, false> > _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _UIntPtrType _M_date_time_formats __iterator_category<char const*> use_facet<std::moneypunct<char, true> > _M_neg_format _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Em __intl __ctr time_get_byname<char, std::istreambuf_iterator<char, std::char_traits<char> > > __add_unsigned<unsigned int> _ZNK9__gnu_cxx17__normal_iteratorIPcSsEixEl _ZNSt17moneypunct_bynameIcLb0EED0Ev _CharT2 _ZNSt17__timepunct_cacheIcEaSERKS0_ __cs2 __cs3 _ZNSt17__timepunct_cacheIcED2Ev mktime __base _ZNSt5__padIcSt11char_traitsIcEE6_S_padERSt8ios_basecPcPKcll _ZNSt18__moneypunct_cacheIcLb0EED0Ev _ZNSt8messagesIcED0Ev _M_thousands_sep __enable_if<true, short unsigned int> __convert_from_v _M_date_formats _ZSt9has_facetISt5ctypeIcEEbRKSt6locale __tm_gmtoff __cs_size _ZNSt16__numpunct_cacheIcED0Ev _ZNKSt10moneypunctIcLb0EE13negative_signEv _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev equal _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10date_orderEv __lo2 _ZN9__gnu_cxx17__normal_iteratorIPcSsEmmEi __testeof _ZN9__gnu_cxx17__normal_iteratorIPcSsEmmEv _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecb do_truename _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecd _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basece _ZSt9use_facetISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _M_initialize_numpunct _ZNKSt10moneypunctIcLb0EE8groupingEv _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecm __max_exp _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecx _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13do_date_orderEv __found_mantissa moneypunct<char, false> moneypunct_byname<char, false> _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe _ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE5equalERKS2_ _ZNKSt8ios_base9precisionEv _M_time_era_format _ZNKSt7collateIcE10do_compareEPKcS2_S2_S2_ _ZSt9has_facetISt7codecvtIcc9mbstate_tEEbRKSt6locale _ZNSt14codecvt_bynameIcc9mbstate_tEC2EPKcm _ZNSt11__timepunctIcE23_M_initialize_timepunctEPi __use_cache<std::__moneypunct_cache<char, true> > __nmatches _ZNK9__gnu_cxx17__normal_iteratorIPKcSsEdeEv __testt _M_insert_int<long long unsigned int> __tmp _ZNKSt8messagesIcE18_M_convert_to_charERKSs __timepunct<char> _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb1EEES3_S3_RSt8ios_basecRKSs _ZNKSt10moneypunctIcLb1EE16do_decimal_pointEv _S_oend __msgid _ZNSt16__numpunct_cacheIcE8_M_cacheERKSt6locale _M_pos_format ~time_get _ZNKSt11__use_cacheISt16__numpunct_cacheIcEEclERKSt6locale _ZNSt10moneypunctIcLb1EEC2EPSt18__moneypunct_cacheIcLb1EEm __mandatory_sign _ZNSt10moneypunctIcLb1EEC2Em ~money_put __hi _ZNKSt7collateIcE12do_transformEPKcS2_ _M_extract_int<short unsigned int> __i1 bidirectional_iterator_tag ~codecvt_byname __cache_type __tmpyear __sep_pos __one __minlen _ZN9__gnu_cxx13new_allocatorIwE8allocateEmPKv _ZN9__gnu_cxx13new_allocatorIwE9constructEPwRKw nothrow_t _ZN9__gnu_cxx13new_allocatorIwE10deallocateEPwm _ZNSaIcEC2ERKS_ _ZNSaIwEC2ERKS_ _ZN9__gnu_cxx13new_allocatorIwE7destroyEPw _ZNSaIwEC2Ev _ZNK9__gnu_cxx13new_allocatorIwE7addressERKw _ZNSaIcEC2Ev _ZNSaIwED2Ev _ZSt7nothrow _ZNK9__gnu_cxx13new_allocatorIwE8max_sizeEv ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/allocator-inst.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=allocator-inst.lo _ZNSaIcED2Ev new_allocator<wchar_t> _ZNK9__gnu_cxx13new_allocatorIwE7addressERw _ZNKSt5ctypeIcE10do_tolowerEc _ZNKSt5ctypeIcE10do_tolowerEPcPKc _ZNSt10ctype_base5lowerE GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=ctype.lo _ZNKSt5ctypeIcE10do_toupperEPcPKc strtok _M_narrow_init strcoll strerror __builtin_memcmp _ZNSt10ctype_base5digitE _M_narrow_ok _ZNKSt5ctypeIcE2isEPKcS2_Pj classic_table do_tolower _ZNSt10ctype_base5alnumE _ZNSt10ctype_base5punctE _M_table _ZNSt10ctype_base5upperE _M_toupper __to_type _ZNSt5ctypeIcED0Ev _ZNKSt5ctypeIcE7tolowerEPcPKc _M_widen _M_del _M_tolower strxfrm _ZNKSt5ctypeIcE7toupperEPcPKc _ZNKSt5ctypeIcE10do_toupperEc _ZNSt10ctype_base5printE _ZNKSt5ctypeIcE5tableEv _M_widen_ok _ZNSt10ctype_base5spaceE ~ctype ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/ctype.cc _ZNSt5ctypeIcE10table_sizeE _ZNSt5ctypeIcE13classic_tableEv _ZNKSt5ctypeIcE9do_narrowEPKcS2_cPc _ZNKSt5ctypeIcE14_M_narrow_initEv _ZNSt10ctype_base5alphaE _ZNSt5ctypeIcE2idE _ZNSt5ctypeIcED2Ev _M_narrow _M_c_locale_ctype _ZNKSt5ctypeIcE7tolowerEc _ZNSt10ctype_base5cntrlE _ZNSt10ctype_base6xdigitE table_size _ZNKSt5ctypeIcE6narrowEPKcS2_cPc _ZNSt10ctype_base5graphE do_toupper is_open buf_cout_sync _ZN14__gnu_internal7buf_cinE __gend _S_synced_with_stdio __tiestr _ZNSt9basic_iosIcSt11char_traitsIcEE5rdbufEPSt15basic_streambufIcS1_E buf_cin_sync buf_cin buf_cerr __sync stdin _ZNKSt13basic_filebufIcSt11char_traitsIcEE7is_openEv _ZN14__gnu_internal13buf_cerr_syncE buf_cout _ZSt4cerr _ZNSt15basic_streambufIcSt11char_traitsIcEE4setgEPcS3_S3_ __atomic_add_single _ZN14__gnu_internal8buf_cerrE __gnu_internal _ZSt4cout _ZNSt8ios_base4InitC2Ev _ZNSt9basic_iosIcSt11char_traitsIcEE3tieEPSo _ZN14__gnu_internal13buf_cout_syncE _ZN14__gnu_internal12buf_cin_syncE _ZNSt8ios_base15sync_with_stdioEb stdio_filebuf<char, std::char_traits<char> > basic_filebuf<char, std::char_traits<char> > __atomic_add_dispatch setg setp ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/ios_init.cc __gnext _ZNSt8ios_base4InitD2Ev GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=ios_init.lo _ZN14__gnu_internal8buf_coutE _ZNSt15basic_streambufIcSt11char_traitsIcEE4setpEPcS3_ _ZSt4clog stderr __pbeg _ZSt3cin __init sync_with_stdio ~Init stdout buf_cerr_sync _ZN9__gnu_cxx4ropeIcSaIcEE26_S_concat_and_set_balancedEPNS_13_Rope_RopeRepIcS1_EES5_ _S_rounded_up_size _ZN9__gnu_cxx4ropeIcSaIcEE5clearEv _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmmPKcm _ZN9__gnu_cxx4ropeIcSaIcEE6insertEmRKS2_ _ZN9__gnu_cxx13_Rope_RopeRepIcSaIcEE12_M_free_treeEv _Placeholder<26> _ZN9__gnu_cxx4ropeIcSaIcEE6insertEmRKNS_14_Rope_iteratorIcS1_EES6_ _ZN9__gnu_cxx4ropeIcSaIcEE6appendERKS2_ reverse_iterator<__gnu_cxx::_Rope_const_iterator<char, std::allocator<char> > > _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED2Ev __left_len _ZNK9__gnu_cxx14_Rope_rep_baseIcSaIcEE13get_allocatorEv _Placeholder<27> _ZN9__gnu_cxx4ropeIcSaIcEE21_S_add_leaf_to_forestEPNS_13_Rope_RopeRepIcS1_EEPS5_ _ZN9__gnu_cxx20_Rope_char_ref_proxyIcSaIcEEaSERKS2_ _S_flatten _L_allocate _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EEc _ZNSt12__basic_fileIcE7seekoffExSt12_Ios_Seekdir _Placeholder<28> _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmRKS2_ _ZNK9__gnu_cxx10_Rope_baseIcSaIcEE13get_allocatorEv _ZN9__gnu_cxx4ropeIcSaIcEE20_S_new_RopeSubstringEPNS_13_Rope_RopeRepIcS1_EEmmRS1_ _Placeholder<29> _ZN9__gnu_cxx14_Rope_rep_baseIcSaIcEE16_M_get_allocatorEv reverse_iterator<__gnu_cxx::_Rope_iterator<char, std::allocator<char> > > _ZN9__gnu_cxx4ropeIcSaIcEE5eraseERKNS_14_Rope_iteratorIcS1_EE _S_deallocate _S_concat_and_set_balanced _ZN9__gnu_cxx10_Rope_baseIcSaIcEE11_F_allocateEm _ZNK9__gnu_cxx4ropeIcSaIcEE15apply_to_piecesEmmRNS_19_Rope_char_consumerIcEE _ZN9__gnu_cxx20_Rope_char_ref_proxyIcSaIcEEaSEc _L_deallocate _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EEPKc showmanyc _ZN9__gnu_cxx4ropeIcSaIcEE10_S_compareEPKNS_13_Rope_RopeRepIcS1_EES6_ _ZNK9__gnu_cxx4ropeIcSaIcEE2atEm _S_destr_leaf_concat_char_iter _ZN9__gnu_cxx4ropeIcSaIcEE6insertEmmc _S_new_RopeLeaf _Swallow_assign _Data_allocate _ZN9__gnu_cxx4ropeIcSaIcEE6insertERKNS_14_Rope_iteratorIcS1_EEc _ZNK9__gnu_cxx4ropeIcSaIcEE4copyEmmPc _ZN9__gnu_cxx4ropeIcSaIcEE5beginEv _ZN9__gnu_cxx14_Rope_RopeLeafIcSaIcEE18_S_rounded_up_sizeEm _ZN9__gnu_cxx14_Rope_rep_baseIcSaIcEE16_Data_deallocateEPcm _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmPKc _ZNKSt12__basic_fileIcE7is_openEv _ZN9__gnu_cxx4ropeIcSaIcEE6insertERKNS_14_Rope_iteratorIcS1_EERKNS_20_Rope_const_iteratorIcS1_EESA_ _ZN9__gnu_cxx4ropeIcSaIcEE9pop_frontEv _ZN9__gnu_cxx4ropeIcSaIcEE6insertERKNS_14_Rope_iteratorIcS1_EEPKcm _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EES6_RKNS_20_Rope_const_iteratorIcS1_EESA_ _S_add_to_forest _ZN9__gnu_cxx13_Rope_RopeRepIcSaIcEE15_M_unref_nonnilEv _ZN9__gnu_cxx4ropeIcSaIcEE19_S_concat_char_iterEPNS_13_Rope_RopeRepIcS1_EEPKcm _M_get_allocator _ZNK9__gnu_cxx4ropeIcSaIcEE6rbeginEv _ZN9__gnu_cxx4ropeIcSaIcEE10push_frontEc _ZN9__gnu_cxx4ropeIcSaIcEE6insertEmRKNS_20_Rope_const_iteratorIcS1_EES6_ _ZN9__gnu_cxx13_Rope_RopeRepIcSaIcEE6_S_refEPS2_ _S_is_roughly_balanced __gthread_mutex_t _S_fetch_ptr _ZN9__gnu_cxx4ropeIcSaIcEE10_S_flattenEPNS_13_Rope_RopeRepIcS1_EEmmPc _S_allocated_capacity _ZN9__gnu_cxx4ropeIcSaIcEE6appendENS_20_Rope_const_iteratorIcS1_EES4_ _ZN9__gnu_cxx10_Rope_baseIcSaIcEE11_C_allocateEm _ZN9__gnu_cxx4ropeIcSaIcEE8pop_backEv _S_dump __filebuf_type _ZN9__gnu_cxx4ropeIcSaIcEE6substrENS_20_Rope_const_iteratorIcS1_EE _M_delete_when_done _M_current_valid _ZNSt12__basic_fileIcE5closeEv _ZNK9__gnu_cxx4ropeIcSaIcEE6substrENS_20_Rope_const_iteratorIcS1_EES4_ _Rope_RopeLeaf<char, std::allocator<char> > _S_is_almost_balanced _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE2fdEv _ZN9__gnu_cxx4ropeIcSaIcEEaSERKS2_ _RC_t _ZN9__gnu_cxx14_Rope_rep_baseIcSaIcEE11_F_allocateEm ~_Rope_RopeFunction _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmPKcS4_ _ZN9__gnu_cxx4ropeIcSaIcEE6insertERKNS_14_Rope_iteratorIcS1_EEmc _ZN9__gnu_cxx4ropeIcSaIcEE6rbeginEv _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EEPKcm _ZN9__gnu_cxx10_Rope_baseIcSaIcEE13_C_deallocateEPNS_23_Rope_RopeConcatenationIcS1_EEm _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EENS_20_Rope_const_iteratorIcS1_EES8_ sys_open _ZN9__gnu_cxx4ropeIcSaIcEE6appendEPKcm _ZNK9__gnu_cxx4ropeIcSaIcEE4findEcm _ZN9__gnu_cxx4ropeIcSaIcEE10_S_balanceEPNS_13_Rope_RopeRepIcS1_EE _Rope_char_ref_proxy _ZN9__gnu_cxx14_Rope_rep_baseIcSaIcEE13_S_deallocateEPNS_19_Rope_RopeSubstringIcS1_EEm ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/ext-inst.cc _ZNSt12__basic_fileIcE4openEPKcSt13_Ios_Openmodei _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EES6_RKS2_ _S_substring _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmmRKNS_20_Rope_const_iteratorIcS1_EES6_ _ZN9__gnu_cxx10_Rope_baseIcSaIcEE11_S_allocateEm _ZN9__gnu_cxx4ropeIcSaIcEE12mutable_rendEv _Data_deallocate const_end mutable_begin _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmPKcm _ZN9__gnu_cxx10_Rope_baseIcSaIcEE11_L_allocateEm _ZNK9__gnu_cxx14_Rope_rep_baseIcSaIcEE16_M_get_allocatorEv _S_allocate _S_leaf _F_deallocate _ZN9__gnu_cxx4ropeIcSaIcEE10_S_flattenEPNS_13_Rope_RopeRepIcS1_EEPc _ZN9__gnu_cxx4ropeIcSaIcEE7balanceEv _S_is_balanced ~rope _ZN9__gnu_cxx18_Rope_RopeFunctionIcSaIcEEaSERKS2_ _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmmPKcS4_ _ZN9__gnu_cxx4ropeIcSaIcEE6insertEmPKcS4_ _ZNSt12__basic_fileIcE8sys_openEP4FILESt13_Ios_Openmode _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmmPKc _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EES6_S6_S6_ _M_free_c_string _ZN9__gnu_cxx4ropeIcSaIcEE12_S_fetch_ptrEPNS_13_Rope_RopeRepIcS1_EEm mutable_rend push_front _Rope_const_iterator<char, std::allocator<char> > _F_allocate _ZNSt13basic_filebufIcSt11char_traitsIcEE5closeEv _M_c_string_lock _S_new_RopeSubstring _ZN9__gnu_cxx4ropeIcSaIcEE24_S_new_RopeConcatenationEPNS_13_Rope_RopeRepIcS1_EES5_RS1_ _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmmc _M_free_tree _ZN9__gnu_cxx4ropeIcSaIcEE18replace_with_c_strEv _ZN9__gnu_cxx14_Rope_rep_baseIcSaIcEE14_Data_allocateEm _ZN9__gnu_cxx13_Rope_RopeRepIcSaIcEE14_S_free_stringEPcmRS1_ _Rope_RopeSubstring<char, std::allocator<char> > _M_cfile_created _M_ref_count _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EES6_PKc const_begin _ZN9__gnu_cxx4ropeIcSaIcEE20mutable_reference_atEm _ZN9__gnu_cxx4ropeIcSaIcEE6insertEm _ZN9__gnu_cxx4ropeIcSaIcEE4dumpEv _Rope_char_consumer<char> _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmc _S_balance _ZN9__gnu_cxx4ropeIcSaIcEE14mutable_rbeginEv _ZN9__gnu_cxx14_Rope_rep_baseIcSaIcEE11_L_allocateEm _S_ref _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EERKS2_ __detail _ZN9__gnu_cxx4ropeIcSaIcEE6_S_refEPNS_13_Rope_RopeRepIcS1_EE _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE4fileEv _Rope_RopeRep<char, std::allocator<char> > _M_depth _ZN9__gnu_cxx4ropeIcSaIcEE12delete_c_strEv pop_back _ZNK9__gnu_cxx4ropeIcSaIcEE10const_rendEv _ZN9__gnu_cxx14_Refcount_Base7_M_decrEv _ZN9__gnu_cxx4ropeIcSaIcEE14_S_is_balancedEPNS_13_Rope_RopeRepIcS1_EE _Refcount_Base _S_min_len __cstr _ZN9__gnu_cxx4ropeIcSaIcEE30_S_destr_leaf_concat_char_iterEPNS_14_Rope_RopeLeafIcS1_EEPKcm _ZN9__gnu_cxx4ropeIcSaIcEE5eraseEmm _ZN9__gnu_cxx4ropeIcSaIcEE15_S_char_ptr_lenEPKc char_producer<char> _ZN9__gnu_cxx4ropeIcSaIcEE9push_backEc _ZN9__gnu_cxx4ropeIcSaIcEE25_S_destr_concat_char_iterEPNS_13_Rope_RopeRepIcS1_EEPKcm _ZN9__gnu_cxx4ropeIcSaIcEE21_S_allocated_capacityEm _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EES6_PKcS8_ _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EEPKcS8_ _S_RopeLeaf_from_unowned_char_ptr mutable_end _ZNK9__gnu_cxx4ropeIcSaIcEEixEm _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2Ev _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmRKNS_14_Rope_iteratorIcS1_EES6_ _S_apply_to_pieces _Placeholder<1> _M_pos _ZN9__gnu_cxx4ropeIcSaIcEE10_S_min_lenE _S_tree_concat _ZN9__gnu_cxx10_Rope_baseIcSaIcEE16_Data_deallocateEPcm _Num _ZN9__gnu_cxx10_Rope_baseIcSaIcEEaSERKS2_ _Placeholder<2> _My_rope _ZN9__gnu_cxx4ropeIcSaIcEE6insertEmc _ZNSt12__basic_fileIcE9showmanycEv _ZN9__gnu_cxx10_Rope_baseIcSaIcEE13_S_deallocateEPNS_19_Rope_RopeSubstringIcS1_EEm delete_c_str _Placeholder<3> _S_concat _ZN9__gnu_cxx14_Rope_rep_baseIcSaIcEE13_F_deallocateEPNS_18_Rope_RopeFunctionIcS1_EEm _ZN9__gnu_cxx10_Rope_baseIcSaIcEE13_L_deallocateEPNS_14_Rope_RopeLeafIcS1_EEm _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EES6_c _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2EiSt13_Ios_Openmodem __basic_file<char> _ZN9__gnu_cxx4ropeIcSaIcEE16_S_add_to_forestEPNS_13_Rope_RopeRepIcS1_EEPS5_ _ZN9__gnu_cxx4ropeIcSaIcEE6insertERKNS_14_Rope_iteratorIcS1_EE _ZN9__gnu_cxx14_Rope_rep_baseIcSaIcEE11_S_allocateEm _ZN9__gnu_cxx4ropeIcSaIcEE11mutable_endEv _Rope_rep_base _Placeholder<4> _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmmRKNS_14_Rope_iteratorIcS1_EES6_ _ZN9__gnu_cxx4ropeIcSaIcEE18_S_rounded_up_sizeEm _M_left mutable_rbegin _ZNK9__gnu_cxx10_Rope_baseIcSaIcEE16_M_get_allocatorEv _Placeholder<5> _M_root _ZN9__gnu_cxx4ropeIcSaIcEE19_S_new_RopeFunctionEPNS_13char_producerIcEEmbRS1_ _ZN9__gnu_cxx13_Rope_RopeRepIcSaIcEEaSERKS2_ _M_set_buffer _ZNSt12__basic_fileIcE8sys_openEiSt13_Ios_Openmode _Placeholder<6> _ZNK9__gnu_cxx4ropeIcSaIcEE11const_beginEv _ZN9__gnu_cxx4ropeIcSaIcEE6insertEmPKc _ZNK9__gnu_cxx4ropeIcSaIcEE9const_endEv _M_fn _ZNK9__gnu_cxx4ropeIcSaIcEE6substrEmm placeholders _Placeholder<7> _M_ref_nonnil _ZNSt13basic_filebufIcSt11char_traitsIcEE13_M_set_bufferEl _ZN9__gnu_cxx4ropeIcSaIcEE33_S_RopeLeaf_from_unowned_char_ptrEPKcmRS1_ _Rope_char_ptr_proxy<char, std::allocator<char> > _ZN9__gnu_cxx4ropeIcSaIcEE22_S_is_roughly_balancedEPNS_13_Rope_RopeRepIcS1_EE _Rope_RopeConcatenation<char, std::allocator<char> > _ZN9__gnu_cxx13_Rope_RopeRepIcSaIcEE16_S_free_if_unrefEPS2_ _ZN9__gnu_cxx14_Refcount_Base7_M_incrEv _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmRKNS_20_Rope_const_iteratorIcS1_EES6_ _S_concat_char_iter _Placeholder<8> operator char _S_add_leaf_to_forest _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2EP4FILESt13_Ios_Openmodem _ZNSt12__basic_fileIcE4fileEv _Rope_base<char, std::allocator<char> > _Rope_iterator<char, std::allocator<char> > _Placeholder<9> __testout _ZNK9__gnu_cxx4ropeIcSaIcEE5frontEv xsputn_2 _M_size _M_decr _M_tag _ZNK9__gnu_cxx4ropeIcSaIcEE8max_sizeEv _M_right _ZN9__gnu_cxx10_Rope_baseIcSaIcEE13_F_deallocateEPNS_18_Rope_RopeFunctionIcS1_EEm _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EES4_S4_ _S_new_RopeConcatenation _M_is_balanced _ZN9__gnu_cxx4ropeIcSaIcEE4rendEv pop_front _ZN9__gnu_cxx14_Rope_rep_baseIcSaIcEE13_C_deallocateEPNS_23_Rope_RopeConcatenationIcS1_EEm _Rope_rep_base<char, std::allocator<char> > _ZN9__gnu_cxx4ropeIcSaIcEE9_S_concatEPNS_13_Rope_RopeRepIcS1_EES5_ _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEPNS_13_Rope_RopeRepIcS1_EEmmS5_ ~basic_filebuf _M_c_string _ZNK9__gnu_cxx4ropeIcSaIcEE4rendEv _ZNK9__gnu_cxx4ropeIcSaIcEE5beginEv _Rope_char_ref_proxy<char, std::allocator<char> > _ZNK9__gnu_cxx4ropeIcSaIcEE12const_rbeginEv _ZN9__gnu_cxx10_Rope_baseIcSaIcEE14_Data_allocateEm __testin _ZNK9__gnu_cxx4ropeIcSaIcEE5emptyEv replace_with_c_str _ZN9__gnu_cxx4ropeIcSaIcEE15_S_new_RopeLeafEPcmRS1_ _ZN9__gnu_cxx4ropeIcSaIcEE7replaceEmmRKS2_ _M_ref_count_lock _ZN9__gnu_cxx4ropeIcSaIcEE6insertERKNS_14_Rope_iteratorIcS1_EES6_S6_ _ZN9__gnu_cxx4ropeIcSaIcEE3endEv _S_unref _ZN9__gnu_cxx4ropeIcSaIcEE13mutable_beginEv _Rope_RopeRep _S_is0 const_rbegin mutable_reference_at _ZNSt13basic_filebufIcSt11char_traitsIcEE27_M_allocate_internal_bufferEv _ZN9__gnu_cxx4ropeIcSaIcEE6appendEc _Tag _ZN9__gnu_cxx4ropeIcSaIcEE4swapERS2_ _ZN9__gnu_cxx4ropeIcSaIcEE6appendEv _ZN9__gnu_cxx4ropeIcSaIcEE7replaceERKNS_14_Rope_iteratorIcS1_EES6_PKcm _Placeholder<10> ~_Rope_RopeLeaf _ZN9__gnu_cxx4ropeIcSaIcEE7_S_dumpEPNS_13_Rope_RopeRepIcS1_EEi _ZNK9__gnu_cxx4ropeIcSaIcEE6substrENS_14_Rope_iteratorIcS1_EE _ZN9__gnu_cxx4ropeIcSaIcEE6insertERKNS_14_Rope_iteratorIcS1_EEPKc _M_cfile _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED0Ev _ZNK9__gnu_cxx4ropeIcSaIcEE6substrENS_14_Rope_iteratorIcS1_EES4_ _ZN9__gnu_cxx4ropeIcSaIcEE6insertEmPKcm _ZN9__gnu_cxx4ropeIcSaIcEE6appendEPKcS4_ _Placeholder<11> _ZSt20__throw_length_errorPKc _ZN9__gnu_cxx4ropeIcSaIcEE5eraseEm _ZN9__gnu_cxx4ropeIcSaIcEE8_S_unrefEPNS_13_Rope_RopeRepIcS1_EE _ZN9__gnu_cxx13_Rope_RopeRepIcSaIcEE13_M_ref_nonnilEv GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=ext-inst.lo _Placeholder<12> _ZNK9__gnu_cxx4ropeIcSaIcEE3endEv _ZNK9__gnu_cxx4ropeIcSaIcEE4copyEPc const_rend _ZNSt12__basic_fileIcE8xsputn_2EPKclS2_l _ZNK9__gnu_cxx4ropeIcSaIcEE4findEPKcm _M_tree_ptr _ZN9__gnu_cxx4ropeIcSaIcEE6appendEPKc _ZNK9__gnu_cxx4ropeIcSaIcEE5c_strEv _S_destr_concat_char_iter _S_free_string _S_substringfn _Placeholder<13> _ZN9__gnu_cxx4ropeIcSaIcEE18_S_apply_to_piecesERNS_19_Rope_char_consumerIcEEPKNS_13_Rope_RopeRepIcS1_EEmm _ZNK9__gnu_cxx4ropeIcSaIcEE4sizeEv ~_Rope_RopeConcatenation _ZNSt12__basic_fileIcE6xsputnEPKcl _S_function _ZN9__gnu_cxx23_Rope_RopeConcatenationIcSaIcEEaSERKS2_ _S_leaf_concat_char_iter _Placeholder<14> _Rope_base _ZN9__gnu_cxx14_Rope_rep_baseIcSaIcEE11_C_allocateEm _ZN9__gnu_cxx14_Rope_rep_baseIcSaIcEE13_L_deallocateEPNS_14_Rope_RopeLeafIcS1_EEm _M_unref_nonnil _ZN9__gnu_cxx4ropeIcSaIcEE6appendEmc _Placeholder<15> ~__basic_file _ZN9__gnu_cxx13_Rope_RopeRepIcSaIcEE8_S_unrefEPS2_ _ZNK9__gnu_cxx4ropeIcSaIcEE4backEv _Placeholder<20> _ZN9__gnu_cxx4ropeIcSaIcEE12_S_substringEPNS_13_Rope_RopeRepIcS1_EEmm _S_fetch _Placeholder<16> _ZN9__gnu_cxx4ropeIcSaIcEE24_S_leaf_concat_char_iterEPNS_14_Rope_RopeLeafIcS1_EEPKcm _ZN9__gnu_cxx4ropeIcSaIcEE8_S_fetchEPNS_13_Rope_RopeRepIcS1_EEm _ZN9__gnu_cxx14_Rope_RopeLeafIcSaIcEEaSERKS2_ _Placeholder<21> _Placeholder<17> _ZN9__gnu_cxx4ropeIcSaIcEE6insertERKNS_14_Rope_iteratorIcS1_EEPKcS8_ _S_new_RopeFunction _S_char_ptr_len _Rope_RopeFunction<char, std::allocator<char> > _ZNSt12__basic_fileIcE2fdEv _C_allocate _Placeholder<22> _ZNK9__gnu_cxx20_Rope_char_ref_proxyIcSaIcEEcvcEv _Placeholder<18> _M_allocate_internal_buffer _ZN9__gnu_cxx4ropeIcSaIcEE5eraseERKNS_14_Rope_iteratorIcS1_EES6_ __fd _S_free_if_unref _ZNK9__gnu_cxx4ropeIcSaIcEE6lengthEv ~stdio_filebuf _ZNSt12__basic_fileIcE4syncEv _Placeholder<23> _ZNK9__gnu_cxx20_Rope_char_ref_proxyIcSaIcEEadEv _Placeholder<19> _ZN9__gnu_cxx4ropeIcSaIcEE6_S_is0Ec _ZN9__gnu_cxx4ropeIcSaIcEE21_S_is_almost_balancedEPNS_13_Rope_RopeRepIcS1_EE __throw_length_error _Placeholder<24> _ZN9__gnu_cxx4ropeIcSaIcEE14_S_tree_concatEPNS_13_Rope_RopeRepIcS1_EES5_ _M_incr _S_empty_c_str _ZN9__gnu_cxx13_Rope_RopeRepIcSaIcEE16_M_free_c_stringEv _ZNK9__gnu_cxx4ropeIcSaIcEE7compareERKS2_ rope<char, std::allocator<char> > __c_lock _ZN9__gnu_cxx4ropeIcSaIcEE6insertERKNS_14_Rope_iteratorIcS1_EERKS2_ _ZNSt12__basic_fileIcE6xsgetnEPcl _C_deallocate _ZN9__gnu_cxx10_Rope_baseIcSaIcEE16_M_get_allocatorEv _Placeholder<25> __wrote ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/streambuf.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=streambuf.lo _M_stringbuf_init _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE17_M_stringbuf_initESt13_Ios_Openmode _M_sync pbase _ZNKSt19basic_ostringstreamIcSt11char_traitsIcESaIcEE3strEv _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEEC1ERKSsSt13_Ios_Openmode _M_string ~basic_stringbuf __capacity __conv _ZNKSt18basic_stringstreamIcSt11char_traitsIcESaIcEE5rdbufEv _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEEC1ESt13_Ios_Openmode __max_size _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEED2Ev _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEED1Ev __newoffo _ZNKSt15basic_streambufIcSt11char_traitsIcEE5pbaseEv _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEEC1ERKSsSt13_Ios_Openmode GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=sstream-inst.lo eback _M_stringbuf basic_istringstream<char, std::char_traits<char>, std::allocator<char> > _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEE3strERKSs _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE3strERKSs __testpos _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEE3strERKSs _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE9underflowEv _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE7seekposESt4fposI9mbstate_tESt13_Ios_Openmode _M_pbump _ZNKSt18basic_stringstreamIcSt11char_traitsIcESaIcEE3strEv _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE15_M_update_egptrEv basic_ostringstream<char, std::char_traits<char>, std::allocator<char> > _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEED0Ev _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEEC2ESt13_Ios_Openmode _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE8_M_pbumpEPcS4_x _ZNKSt15basic_stringbufIcSt11char_traitsIcESaIcEE3strEv _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE9pbackfailEi _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE6setbufEPcl _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE7_M_syncEPcmm _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEEC2ERKSsSt13_Ios_Openmode _ZNKSt15basic_streambufIcSt11char_traitsIcEE5ebackEv __testput _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEEC2ERKSsSt13_Ios_Openmode __string_type _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEED0Ev __endp __testeq _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEEC2ESt13_Ios_Openmode _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEEC1ESt13_Ios_Openmode basic_iostream<char, std::char_traits<char> > _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEED1Ev _ZNSs12_S_constructIPcEES0_T_S1_RKSaIcESt20forward_iterator_tag ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/sstream-inst.cc _ZNSs12_S_constructIPcEES0_T_S1_RKSaIcE ~basic_stringstream __is_null_pointer<char> basic_stringstream<char, std::char_traits<char>, std::allocator<char> > _M_mode __endg __distance<char*> __newoffi ~basic_ostringstream ~basic_istream max<long unsigned int> _ZNKSt19basic_istringstreamIcSt11char_traitsIcESaIcEE3strEv _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEED2Ev _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEED2Ev _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEE3strERKSs __stringbuf_type _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE9showmanycEv _ZNKSt19basic_ostringstreamIcSt11char_traitsIcESaIcEE5rdbufEv _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEEC2ESt13_Ios_Openmode _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEEC1ERKSsSt13_Ios_Openmode _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE8overflowEi __testboth _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEED0Ev _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEED1Ev _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEEC1ESt13_Ios_Openmode _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEED0Ev _S_construct_aux<char*> _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEEC2ESt13_Ios_Openmode _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEEC2ERKSsSt13_Ios_Openmode _S_construct<char*> _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEEC2ERKSsSt13_Ios_Openmode __iterator_category<char*> ~basic_iostream basic_string<char*> _M_update_egptr __opt_len ~basic_istringstream _ZNKSt19basic_istringstreamIcSt11char_traitsIcESaIcEE5rdbufEv _ZNSs16_S_construct_auxIPcEES0_T_S1_RKSaIcESt12__false_type basic_stringbuf<char, std::char_traits<char>, std::allocator<char> > _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEED2Ev is_bounded _ZNSt8ios_base6eofbitE _M_iword _ZNSt8ios_base3decE is_specialized _M_streambuf_state _ZNSt8ios_base8internalE has_infinity _ZNSt8ios_base9boolalphaE has_denorm _ZNSt8ios_base6binaryE is_iec559 _ZNSt8ios_base5imbueERKSt6locale _ZNSt8ios_base10floatfieldE _ZNSt14numeric_limitsIiE3maxEv _ZNSt8ios_base7_M_initEv _ZNSt8ios_base6skipwsE _ZNSt8ios_base4leftE _S_top _M_ios_locale _M_call_callbacks is_exact ~ios_base _ZNSt8ios_base14_Callback_list19_M_remove_referenceEv _ZNSt8ios_base8showbaseE _ZNSt8ios_base6xallocEv _ZNSt8ios_base2inE _M_word _ZNSt8ios_base4Init20_S_synced_with_stdioE _M_word_size _ZNSt8ios_base20_M_dispose_callbacksEv event_callback _ZNSt14numeric_limitsIiE9quiet_NaNEv xalloc _ZNSt8ios_base7goodbitE _M_exception digits10 _ZNSt14numeric_limitsIiE11round_errorEv _ZNSt8ios_base3hexE _ZNSt8ios_base3octE is_integer _M_dispose_callbacks denorm_indeterminate ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/ios.cc _ZNSt8ios_baseC2Ev denorm_absent _ZNSt8ios_base4Init11_S_refcountE _ZNSt8ios_base5fixedE _ZNSt8ios_base11adjustfieldE _M_precision _ZSt19__throw_ios_failurePKc max_exponent10 _ZNSt8ios_base9basefieldE _ZNSt8ios_base9showpointE numeric_limits<int> _ZNSt8ios_base6badbitE unsetf imbue_event _ZNSt8ios_base3ateE float_round_style _ZNSt8ios_base10scientificE _ZNSt8ios_base5pwordEi _S_local_word_size _ZNSt8ios_base17register_callbackEPFvNS_5eventERS_iEi _ZNSt8ios_base5truncE _ZNSt8ios_baseaSERKS_ round_indeterminate max_exponent _ZNSt14numeric_limitsIiE10denorm_minEv has_quiet_NaN __cb round_to_nearest round_toward_zero _M_local_word _ZNSt8ios_baseD2Ev _ZNSt8ios_base6unsetfESt13_Ios_Fmtflags _ZNSt14numeric_limitsIiE7epsilonEv __newsize float_denorm_style has_signaling_NaN _ZNSt8ios_base5rightE is_modulo _ZNSt8ios_base14_Callback_list16_M_add_referenceEv _ZNSt14numeric_limitsIiE8infinityEv round_toward_infinity _ZNSt8ios_base9uppercaseE _M_callbacks __words _ZNSt8ios_base17_M_call_callbacksENS_5eventE register_callback _M_init _ZNSt14numeric_limitsIiE3minEv _Callback_list erase_event tinyness_before __iword round_toward_neg_infinity is_signed _ZNSt14numeric_limitsIiE13signaling_NaNEv __next _ZNSt8ios_base3begE _ZNSt8ios_base3appE _M_word_zero __fn __ix epsilon _vptr.ios_base _M_flags __throw_ios_failure _ZNSt8ios_base5iwordEi _ZNSt8ios_base3outE denorm_min _Words traps _ZNSt8ios_base7unitbufE min_exponent denorm_present _ZNSt8ios_base7failbitE has_denorm_loss _M_next round_error __index copyfmt_event _M_grow_words radix _ZNSt8ios_base7showposE _ZNSt8ios_baseD0Ev _ZNSt8ios_base3curE _ZNSt8ios_base3endE GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=ios.lo _M_pword _ZNSt8ios_base13_M_grow_wordsEib _M_width min_exponent10 _ZNSt10__num_base11_S_atoms_inE _ZNSt10money_base8_S_atomsE __fptr __fltfield _ZNSt10money_base18_S_default_patternE GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=locale_facets.lo ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/locale_facets.cc __test _ZNSt17__timepunct_cacheIcE12_S_timezonesE _ZNSt10__num_base12_S_atoms_outE _S_c_locale ~__scoped_lock __newf __cat _S_c_name __is_char<char> __new_size __idpp __fpr _ZNSt6locale4noneE _ZNSt6localeC2EPNS_5_ImplE _ZNKSt6locale5facet19_M_remove_referenceEv _ZN9__gnu_cxx7__mutex6unlockEv _S_single __throw_runtime_error _ZNSt6locale5ctypeE _ZNSt6locale5_ImplC2ERKS0_m _ZNSt6locale5facet18_S_initialize_onceEv _ZNSt6locale10_S_classicE gthread_mutex _ZNSt6locale7numericE _M_device _ZNSt6locale2id11_S_refcountE _ZNSt6locale7collateE _ZNSt6locale8messagesE __oldc __oldf GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=locale.lo __idp _ZNSt6locale5_ImplD2Ev _ZN9__gnu_cxx7__mutex4lockEv _ZNSt6locale5facet11_S_c_localeE _ZN9__gnu_cxx7__mutex13gthread_mutexEv _ZNSt6locale5facetD2Ev _Lock_policy get_locale_cache_mutex _S_atomic _ZNSt6localeC2ERKS_ _ZNKSt6locale5facet16_M_add_referenceEv __enable_if<true, bool> __cpr _ZNSt6locale5facet20_S_lc_ctype_c_localeEPiPKc _S_mutex __newc __fp __mutex _S_categories_size _vptr.facet __imp _ZSt21__throw_runtime_errorPKc _ZNSt6locale8monetaryE __cxa_guard_release __ip __mutex_type ~facet _ZNSt6locale9_S_globalE _ZN9__gnu_cxx13__scoped_lockaSERKS0_ __other _ZNSt6locale5facet9_S_c_nameE _S_lc_ctype_c_locale _ZNSt6locale3allE _ZNSt6locale5facetaSERKS0_ ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/locale.cc __cxa_guard_acquire _ZNSt6locale4timeE _ZNSt6locale5facetD0Ev _ZN9__gnu_cxx7__mutexaSERKS0_ _ZNSt6localeD2Ev _M_mutex __default_lock_policy pubimbue __remaining _ZNSt15basic_streambufIcSt11char_traitsIcEE7seekposESt4fposI9mbstate_tESt13_Ios_Openmode _M_out_end sputbackc _ZNSt15basic_streambufIcSt11char_traitsIcEE8in_availEv _ZNSt15basic_streambufIcSt11char_traitsIcEEC2Ev _ZSt17__copy_streambufsIcSt11char_traitsIcEElPSt15basic_streambufIT_T0_ES6_ _ZNSt15basic_streambufIcSt11char_traitsIcEE7sungetcEv _M_buf_locale _ZNSt15basic_streambufIcSt11char_traitsIcEE8overflowEi _ZNSt15basic_streambufIcSt11char_traitsIcEE9showmanycEv _M_out_beg stossc _ZNSt15basic_streambufIcSt11char_traitsIcEED2Ev _ZNSt15basic_streambufIcSt11char_traitsIcEE9pubsetbufEPcl pubsetbuf _ZNSt15basic_streambufIcSt11char_traitsIcEE6xsputnEPKcl _ZNSt15basic_streambufIcSt11char_traitsIcEEC2ERKS2_ _ZNSt15basic_streambufIcSt11char_traitsIcEE5uflowEv GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=streambuf-inst.lo _M_in_cur _ZNSt15basic_streambufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZNSt15basic_streambufIcSt11char_traitsIcEE6xsgetnEPcl ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/streambuf-inst.cc _ZNSt15basic_streambufIcSt11char_traitsIcEE9pbackfailEi _M_in_end _ZNSt15basic_streambufIcSt11char_traitsIcEE9sputbackcEc _vptr.basic_streambuf _ZNSt15basic_streambufIcSt11char_traitsIcEE5imbueERKSt6locale _M_in_beg _ZNSt15basic_streambufIcSt11char_traitsIcEED0Ev _ZNSt15basic_streambufIcSt11char_traitsIcEE12__safe_pbumpEl _ZNKSt15basic_streambufIcSt11char_traitsIcEE6getlocEv _ZNSt15basic_streambufIcSt11char_traitsIcEE9underflowEv __safe_pbump _ZNSt15basic_streambufIcSt11char_traitsIcEE8pubimbueERKSt6locale _ZNSt15basic_streambufIcSt11char_traitsIcEE5sgetnEPcl _ZNSt15basic_streambufIcSt11char_traitsIcEE6setbufEPcl __buf_len in_avail _M_out_cur sungetc _ZNSt15basic_streambufIcSt11char_traitsIcEE4syncEv _ZNSt15basic_streambufIcSt11char_traitsIcEE6stosscEv _ZNSt15basic_streambufIcSt11char_traitsIcEEaSERKS2_ _ZNSt9basic_iosIcSt11char_traitsIcEE15_M_cache_localeERKSt6locale _ZNSt9basic_iosIcSt11char_traitsIcEE7copyfmtERKS2_ __num_get_type __except _ZNKSt9basic_iosIcSt11char_traitsIcEE6narrowEcc _M_fill operator! _M_num_get copyfmt operator void* _M_fill_init _ZNSt9basic_iosIcSt11char_traitsIcEED0Ev _M_ctype _ZNSt9basic_iosIcSt11char_traitsIcEEC2Ev ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/ios-inst.cc _ZNSt9basic_iosIcSt11char_traitsIcEEC2EPSt15basic_streambufIcS1_E GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=ios-inst.lo _M_cache_locale _M_streambuf _M_num_put _ZNKSt9basic_iosIcSt11char_traitsIcEE3badEv _ZNKSt9basic_iosIcSt11char_traitsIcEE3eofEv _ZNSt9basic_iosIcSt11char_traitsIcEED2Ev _ZNSt9basic_iosIcSt11char_traitsIcEE5imbueERKSt6locale _ZNSt9basic_iosIcSt11char_traitsIcEE10exceptionsESt12_Ios_Iostate _M_tie _ZNKSt9basic_iosIcSt11char_traitsIcEEntEv _ZNKSt9basic_iosIcSt11char_traitsIcEEcvPvEv do_encoding __codecvt_abstract_base<char, char, mbstate_t> _ZNSt7codecvtIcc9mbstate_tEC2EPim _ZNSt7codecvtIcc9mbstate_tE2idE _ZNSt7codecvtIcc9mbstate_tED2Ev _ZNKSt7codecvtIcc9mbstate_tE9do_lengthERS0_PKcS4_m GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=codecvt.lo do_out ~__codecvt_abstract_base do_unshift do_length _ZNKSt7codecvtIcc9mbstate_tE10do_unshiftERS0_PcS3_RS3_ __from intern_type __from_next _ZNKSt7codecvtIcc9mbstate_tE11do_encodingEv _ZNKSt7codecvtIcc9mbstate_tE6do_outERS0_PKcS4_RS4_PcS6_RS6_ _ZNKSt7codecvtIcc9mbstate_tE16do_always_noconvEv codecvt_base _M_c_locale_codecvt __to_next partial ~codecvt _ZNSt7codecvtIcc9mbstate_tEC2Em _ZNSt7codecvtIcc9mbstate_tED0Ev _ZNKSt7codecvtIcc9mbstate_tE13do_max_lengthEv do_in extern_type do_max_length _ZNKSt7codecvtIcc9mbstate_tE5do_inERS0_PKcS4_RS4_PcS6_RS6_ ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/codecvt.cc do_always_noconv _ZNSt10moneypunctIcLb1EED0Ev GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=monetary_members.lo monetary_members.cc _ZNSt10moneypunctIcLb0EED2Ev _ZNSt10moneypunctIcLb1EED2Ev _ZNSt10moneypunctIcLb0EED0Ev _ZNSt13basic_filebufIcSt11char_traitsIcEE5imbueERKSt6locale _ZNSt13basic_filebufIcSt11char_traitsIcEED0Ev __computed_off __enc __iresume _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1ERKSsSt13_Ios_Openmode _ZNSt13basic_filebufIcSt11char_traitsIcEE14_M_get_ext_posER9mbstate_t _M_pback _ZNSs5frontEv uint16_t __builtin_memmove _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode _ZNSt13basic_filebufIcSt11char_traitsIcEE4openERKSsSt13_Ios_Openmode _ZNSt14basic_ofstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode _ZNSt14basic_ifstreamIcSt11char_traitsIcEE7is_openEv __blen __avail _ZNSt14basic_ifstreamIcSt11char_traitsIcEE4openERKSsSt13_Ios_Openmode uint_fast32_t _M_codecvt_tmp _ZNKSt23__codecvt_abstract_baseIcc9mbstate_tE8encodingEv _ZNSt13basic_fstreamIcSt11char_traitsIcEE5closeEv _ZNSt13basic_filebufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode __from_end uintmax_t _M_pback_cur_save __file_off _ZNSt13basic_filebufIcSt11char_traitsIcEE19_M_terminate_outputEv _M_seek GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=fstream-inst.lo __ibuf _M_state_cur _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1Ev _ZNSt14basic_ifstreamIcSt11char_traitsIcEE5closeEv _ZNSt14basic_ifstreamIcSt11char_traitsIcEED0Ev _M_pback_init __st _ZNSt13basic_filebufIcSt11char_traitsIcEE15_M_create_pbackEv _M_ext_buf_size piecewise_construct_t _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1ERKSsSt13_Ios_Openmode _ZNSs13shrink_to_fitEv _ZNSt13basic_filebufIcSt11char_traitsIcEE7seekposESt4fposI9mbstate_tESt13_Ios_Openmode _M_ext_next uint_least32_t _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2Ev _M_buf _ZNSt13basic_filebufIcSt11char_traitsIcEE7_M_seekExSt12_Ios_Seekdir9mbstate_t _ZNSt14basic_ifstreamIcSt11char_traitsIcEED1Ev _ZNKSt23__codecvt_abstract_baseIcc9mbstate_tE2inERS0_PKcS4_RS4_PcS6_RS6_ _ZNSt13basic_fstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode _ZZNSt13basic_filebufIcSt11char_traitsIcEE5closeEvEN14__close_sentryD2Ev _ZNSt13basic_fstreamIcSt11char_traitsIcEED1Ev _M_buf_allocated _ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEESt16initializer_listIcE _M_reading basic_ofstream<char, std::char_traits<char> > __bufavail _ZNKSt14basic_ofstreamIcSt11char_traitsIcEE7is_openEv _ZNKSt13basic_fstreamIcSt11char_traitsIcEE7is_openEv _M_buf_size _ZNSt14basic_ifstreamIcSt11char_traitsIcEED2Ev _ZNSt13basic_fstreamIcSt11char_traitsIcEE4openERKSsSt13_Ios_Openmode _ZNSt13basic_filebufIcSt11char_traitsIcEE4syncEv _M_state_last __limit _ZNKSt14basic_ifstreamIcSt11char_traitsIcEE5rdbufEv _ZNKSt23__codecvt_abstract_baseIcc9mbstate_tE10max_lengthEv _M_destroy_internal_buffer _ZNSt13basic_fstreamIcSt11char_traitsIcEEC2ERKSsSt13_Ios_Openmode _ZNKSt14basic_ofstreamIcSt11char_traitsIcEE5rdbufEv uint_least64_t crend _ZNKSs5frontEv _ZNSt13basic_filebufIcSt11char_traitsIcEE26_M_destroy_internal_bufferEv _ZNSt14basic_ofstreamIcSt11char_traitsIcEE5closeEv _ZNSt14basic_ofstreamIcSt11char_traitsIcEE4openERKSsSt13_Ios_Openmode _ZNSt13basic_filebufIcSt11char_traitsIcEE6xsgetnEPcl __got_eof _M_ext_buf _ZNKSt13basic_fstreamIcSt11char_traitsIcEE5rdbufEv _ZNKSt23__codecvt_abstract_baseIcc9mbstate_tE13always_noconvEv piecewise_construct uint_fast16_t _ZNSt13basic_filebufIcSt11char_traitsIcEE9showmanycEv _ZNSt14basic_ofstreamIcSt11char_traitsIcEE7is_openEv _ZNSt13basic_filebufIcSt11char_traitsIcEEC2Ev _ZNSt13basic_filebufIcSt11char_traitsIcEE9underflowEv char32_t _M_lock _ZNSt13basic_fstreamIcSt11char_traitsIcEED0Ev __bend _ZNSs4backEv _ZNSs8pop_backEv _ZNKSs6cbeginEv _ZNSt14basic_ofstreamIcSt11char_traitsIcEED0Ev _ZNSt13basic_filebufIcSt11char_traitsIcEE16_M_destroy_pbackEv _ZNKSt23__codecvt_abstract_baseIcc9mbstate_tE3outERS0_PKcS4_RS4_PcS6_RS6_ cend _ZNKSs7crbeginEv operator!=<mbstate_t> __codecvt_type _ZNSt13basic_fstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode _M_writing _M_ext_end __check_facet<std::codecvt<char, char, mbstate_t> > uintptr_t _ZNSs6appendESt16initializer_listIcE ~basic_fstream cbegin ~basic_ifstream _ZNSt14basic_ofstreamIcSt11char_traitsIcEED1Ev _ZNSt13basic_fstreamIcSt11char_traitsIcEEC1ERKSsSt13_Ios_Openmode uint_least16_t _ZNSt13basic_filebufIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode _ZNSt13basic_filebufIcSt11char_traitsIcEE8overflowEi _M_pback_end_save __remainder __elen _M_destroy_pback _ZNSsaSEOSs _M_terminate_output _M_filebuf uint_fast64_t _ZNKSt23__codecvt_abstract_baseIcc9mbstate_tE7unshiftERS0_PcS3_RS3_ ~__close_sentry __buflen uint_least8_t _ZNSt13basic_filebufIcSt11char_traitsIcEE9pbackfailEi _ZNSt14basic_ofstreamIcSt11char_traitsIcEED2Ev _ZNSspLESt16initializer_listIcE _ZNSt14basic_ifstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode basic_ifstream<char, std::char_traits<char> > _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2ERKSsSt13_Ios_Openmode __rlen _ZNSs6assignESt16initializer_listIcE ~basic_ofstream _ZNKSs4cendEv __buffill _ZNSt13basic_filebufIcSt11char_traitsIcEE6xsputnEPKcl _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_St16initializer_listIcE _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1Ev _M_state_beg __no_movement _ZNSt13basic_fstreamIcSt11char_traitsIcEEC1Ev /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/src/c++11 _M_codecvt _ZNSsaSESt16initializer_listIcE __testpb _M_get_ext_pos __to_end _ZNSt13basic_filebufIcSt11char_traitsIcEE22_M_convert_to_externalEPcl __file_type _ZNSt13basic_fstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode _ZNKSt14basic_ifstreamIcSt11char_traitsIcEE7is_openEv _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2Ev basic_fstream<char, std::char_traits<char> > __gptr_off _ZNSt13basic_fstreamIcSt11char_traitsIcEED2Ev __iend _ZNSt13basic_fstreamIcSt11char_traitsIcEEC2Ev __fbi _ZNKSs4backEv _ZNSt13basic_fstreamIcSt11char_traitsIcEE7is_openEv _ZNKSs5crendEv char16_t shrink_to_fit __fb _M_create_pback _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode _ZNSt13basic_filebufIcSt11char_traitsIcEE6setbufEPcl uint_fast8_t ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11/fstream-inst.cc __chunk initializer_list<char> crbegin _ZNSs6assignEOSs _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2ERKSsSt13_Ios_Openmode __state_type _ZNKSt23__codecvt_abstract_baseIcc9mbstate_tE6lengthERS0_PKcS4_m _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode _M_convert_to_external _ZNSt13basic_filebufIcSt11char_traitsIcEED2Ev __iterator_traits<__gnu_cxx::__normal_iterator<char const*, std::basic_string<char, std::char_traits<char>, std::allocator<char> > >, true> _ZNSsC2IN9__gnu_cxx17__normal_iteratorIPcSsEEEET_S4_RKSaIcE _ZNKSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPKcSsEEEptEv _Tp1 _ZNKSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPKcSsEEEixEl operator+<char, std::char_traits<char>, std::allocator<char> > __osize __n1 __n2 _ZNKSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPcSsEEEmiEl __requested_cap _ZNKSt16initializer_listIcE4sizeEv _ZNSsC2IPcEET_S1_RKSaIcE __req _ZNSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPKcSsEEEmIEl _ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_EPKS3_RKS6_ __is_null_pointer<__gnu_cxx::__normal_iterator<char*, std::basic_string<char> > > _ZNSsC2IPKcEET_S2_RKSaIcE _ZNSsC2ERKSsmmRKSaIcE __distance<__gnu_cxx::__normal_iterator<char*, std::basic_string<char> > > _ZNSs4nposE __malloc_header_size operator-<char const*, std::basic_string<char> > __iterator_traits<__gnu_cxx::__normal_iterator<char*, std::basic_string<char, std::char_traits<char>, std::allocator<char> > >, true> __data rebind<char> _ZNSsC2EPKcmRKSaIcE _ZNSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPcSsEEEmmEi _ZNSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPcSsEEEmmEv _ZNKSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPKcSsEEEplEl _ZNSsC2ERKSs operator!=<char*, std::basic_string<char> > operator==<char const*, std::basic_string<char> > _ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_ERKS6_S8_ _Result _ZNKSt16initializer_listIcE5beginEv __pos1 __pos2 __len1 __len2 _ZNSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPKcSsEEEppEi _ZNKSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPcSsEEEptEv _ZNSs4_Rep20_S_empty_rep_storageE _ZNSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPKcSsEEEppEv _ZNSs12_S_constructIN9__gnu_cxx17__normal_iteratorIPcSsEEEES2_T_S4_RKSaIcESt20forward_iterator_tag _ZNSsC2EPKcRKSaIcE __iterator_category<__gnu_cxx::__normal_iterator<char*, std::basic_string<char> > > iterator<std::random_access_iterator_tag, char, long int, char*, char&> __alloc _ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_ES3_RKS6_ ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11/string-inst.cc _ZNSs12_Alloc_hiderC2EPcRKSaIcE less<char const*> _ZNSsC2Ev __extra _ZNSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPcSsEEEpLEl __throw_logic_error GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=string-inst.lo _S_construct<__gnu_cxx::__normal_iterator<char*, std::basic_string<char> > > _S_construct_aux<__gnu_cxx::__normal_iterator<char*, std::basic_string<char> > > _ZNKSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPcSsEEEdeEv __how_much _ZNKSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPcSsEEEixEl _ZN9__gnu_cxxeqIPKcSsEEbRKNS_17__normal_iteratorIT_T0_EES8_ _ZNSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPKcSsEEEmmEi _ZNSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPKcSsEEEmmEv __adj_size __alloc1 __alloc2 iterator_type _ZNKSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPcSsEEE4baseEv __nleft _ZNSsC2ESt16initializer_listIcERKSaIcE _M_array __pagesize basic_string<__gnu_cxx::__normal_iterator<char*, std::basic_string<char> > > _Arg1 _Arg2 __old_capacity _ZN9__gnu_cxxeqIPcSsEEbRKNS_17__normal_iteratorIT_T0_EES7_ _ZNSs4_Rep11_S_terminalE __old_size _ZNKSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPKcSsEEEmiEl _ZNKSt16initializer_listIcE3endEv _ZSt19__throw_logic_errorPKc _ZNKSt4lessIPKcEclERKS1_S4_ binary_function<char const*, char const*, bool> _ZNKSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPKcSsEEEdeEv __position _ZNKSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPKcSsEEE4baseEv _ZNKSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPcSsEEEplEl _ZNSsC2EmcRKSaIcE _ZNSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPcSsEEEmIEl operator==<char*, std::basic_string<char> > _ZNSs4_Rep11_S_max_sizeE __place _ZNSsC2EOSs _ZNSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPKcSsEEEpLEl iterator<std::random_access_iterator_tag, char, long int, char const*, char const&> initializer_list _ZNSsC2ERKSaIcE _Raw_bytes_alloc _ZNSsD2Ev _ZNSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPcSsEEEppEi _ZNSt16reverse_iteratorIN9__gnu_cxx17__normal_iteratorIPcSsEEEppEv _ZNSsC2ERKSsmm _M_len __gnuc_va_list _ZNKSt15error_condition7messageEv make_error_code _ZSt16generic_categoryv _ZNKSt15error_conditioncvbEv allocator_arg _S_error_space _S_error_stack __throw_overflow_error defer_lock_t _ZNKSt10error_code23default_error_conditionEv _ZNSt10error_code5clearEv _ZNKSt10error_code7messageEv promise_already_satisfied __throw_bad_alloc _M_cat _ZN9__gnu_cxx15__snprintf_liteEPcmPKcS0_ chrono _ZNSt10error_code6assignEiRKSt14error_category __throw_out_of_range __throw_bad_exception _ZSt23__throw_underflow_errorPKc _ZSt19__throw_regex_errorNSt15regex_constants10error_typeE _S_error_badrepeat adopt_lock _ZSt22__throw_overflow_errorPKc ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11/functexcept.cc _ZNSt15error_condition6assignEiRKSt14error_category _ZSt15future_categoryv __throw_underflow_error _ZNKSt15error_condition5valueEv __throw_system_error __throw_regex_error _ZSt17__throw_bad_allocv __throw_future_error _S_error_brace _S_error_brack _S_error_range generic_category _ZNKSt10error_code8categoryEv _ZSt20__throw_system_errori __ap _S_error_paren future_already_retrieved _S_error_collate default_error_condition _ZSt20__throw_domain_errorPKc _ZSt18__throw_bad_typeidv _ZSt25__throw_bad_function_callv _S_error_ctype _S_error_escape __ec _ZNKSt15error_condition8categoryEv _S_error_badbrace _ZNSt15error_condition5clearEv __throw_bad_typeid _M_value __ecode GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=functexcept.lo _ZSt21__throw_bad_exceptionv no_state error_type future_errc try_to_lock __throw_range_error broken_promise defer_lock future_category _ZSt20__throw_out_of_rangePKc _S_error_complexity _ZSt19__throw_range_errorPKc __throw_domain_error allocator_arg_t adopt_lock_t _ZSt24__throw_invalid_argumentPKc _ZSt20__throw_future_errori __throw_bad_function_call _ZNKSt10error_codecvbEv __errc message __snprintf_lite regex_constants __alloca_size try_to_lock_t __throw_invalid_argument _ZNKSt10error_code5valueEv _S_error_backref _ZNSt11regex_errorD0Ev _ZNSt11regex_errorD2Ev ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11/regex.cc _M_code GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=regex.lo ~regex_error _ZNSt11regex_errorC2ENSt15regex_constants10error_typeE _ZNKSt11regex_error4codeEv __istream_type ../../../../gcc-4.9.1/libstdc++-v3/src/c++98/compatibility.cc /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libstdc++-v3/src GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=compatibility.lo _ZNSi6ignoreEv _ZNSt8bad_castD2Ev GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=bad_cast.lo ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/bad_cast.cc what _ZNSt8bad_castD0Ev _ZNKSt8bad_cast4whatEv ~bad_cast _ZN10__cxxabiv121__vmi_class_type_infoD2Ev __virtual_mask __base_info _ZNKSt9type_infoeqERKS_ src_type _ZN10__cxxabiv117__class_type_info16__dyncast_resultaSERKS1_ _ZNK10__cxxabiv121__vmi_class_type_info11__do_upcastEPKNS_17__class_type_infoEPKvRNS1_15__upcast_resultE again contained_p nonvirtual_base_type __is_virtual_p part2dst __offset_flags dst2src _ZNK10__cxxabiv122__base_class_type_info13__is_public_pEv __contained_ambig _ZNK10__cxxabiv117__class_type_info17__find_public_srcElPKvPKS0_S2_ base_access vtable result2_ambig __contained_virtual_mask __contained_mask __do_dyncast new_sub_kind __find_public_src _ZNK10__cxxabiv122__base_class_type_info8__offsetEv __hwm_bit __sub_kind __unknown __public_mask base_kind __upcast_result convert_to_base __contained_private src2dst __base_class_type_info ~__vmi_class_type_info __offset_shift __do_upcast result2 __dyncast_result _ZNK10__cxxabiv122__base_class_type_info14__is_virtual_pEv __do_find_public_src whole2src src_details __arg result_ambig whole2dst __flags_unknown_mask __contained_public_mask dst_cand __base_count old_sub_kind __not_contained _ZN10__cxxabiv121__vmi_class_type_infoD0Ev dst_ptr __diamond_shaped_mask _ZNK10__cxxabiv117__class_type_info11__do_upcastEPKS0_PKvRNS0_15__upcast_resultE ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/vmi_class_type_info.cc __offset_flags_masks is_virtual dst_type obj_ptr _ZNK10__cxxabiv121__vmi_class_type_info20__do_find_public_srcElPKvPKNS_17__class_type_infoES2_ _ZNK10__cxxabiv121__vmi_class_type_info12__do_dyncastElNS_17__class_type_info10__sub_kindEPKS1_PKvS4_S6_RNS1_16__dyncast_resultE details_ __base_type is_public whole_details skip_on_first_pass access_path src_ptr __offset __is_public_p GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=vmi_class_type_info.lo adjust_pointer<void> __flags_masks __non_diamond_repeat_mask __contained_public adjust_pointer<long int> GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=del_opv.lo ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/del_opv.cc ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/eh_globals.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=eh_globals.lo __gxx_caught_object exceptionObject ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/eh_catch.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=eh_catch.lo __cxa_get_exception_ptr _Unwind_DeleteException objectp _ZNKSt9exception4whatEv _ZN10__cxxabiv115__forced_unwind12__pure_dummyEv ~bad_exception _vptr.__forced_unwind ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/eh_exception.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=eh_exception.lo _ZN10__cxxabiv119__foreign_exceptionD2Ev ~__forced_unwind _ZN10__cxxabiv115__forced_unwindD0Ev _ZNSt9exceptionD2Ev _ZNSt13bad_exceptionD2Ev _ZN10__cxxabiv119__foreign_exceptionD0Ev _ZN10__cxxabiv119__foreign_exception12__pure_dummyEv _ZN10__cxxabiv115__forced_unwindD2Ev _ZNSt9exceptionD0Ev _vptr.__foreign_exception ~__foreign_exception __pure_dummy ~exception _ZNKSt13bad_exception4whatEv _vptr.exception _ZNSt13bad_exceptionD0Ev __is_pointer_p ~type_info _ZNKSt9type_info4nameEv _ZNSt9type_infoaSERKS_ _ZNKSt9type_info15__is_function_pEv _vptr.type_info _ZNSt9type_infoD2Ev __do_catch _ZNKSt9type_info11__do_upcastEPKN10__cxxabiv117__class_type_infoEPPv _ZNKSt9type_info14__is_pointer_pEv _ZNKSt9type_info10__do_catchEPKS_PPvj _ZNSt9type_infoD0Ev GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=tinfo.lo __is_function_p thr_type ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/tinfo.cc _ZNKSt9type_info6beforeERKS_ _ZNKSt9type_infoneERKS_ GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=class_type_info.lo _ZNK10__cxxabiv117__class_type_info11__do_upcastEPKS0_PPv ~__class_type_info ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/class_type_info.cc _ZNK10__cxxabiv117__class_type_info10__do_catchEPKSt9type_infoPPvj outer thr_obj _ZN10__cxxabiv117__class_type_infoD0Ev _ZNK10__cxxabiv117__class_type_info12__do_dyncastElNS0_10__sub_kindEPKS0_PKvS3_S5_RNS0_16__dyncast_resultE _ZN10__cxxabiv117__class_type_infoD2Ev contained_public_p _ZN10__cxxabiv117__class_type_infoaSERKS0_ _ZNK10__cxxabiv117__class_type_info20__do_find_public_srcElPKvPKS0_S2_ ~bad_alloc _ZNSt9bad_allocD2Ev _ZNSt9bad_allocD0Ev GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=bad_alloc.lo _ZNKSt9bad_alloc4whatEv ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/bad_alloc.cc __unexpected_handler func _ZSt13set_terminatePFvvE GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=eh_terminate.lo __terminate_handler ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/eh_terminate.cc set_terminate _ZN10__cxxabiv120__unexpected_handlerE set_unexpected _ZSt14set_unexpectedPFvvE _ZN10__cxxabiv119__terminate_handlerE __cxa_guard_abort GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=guard.lo __guard throw_recursive_init_exception set_init_in_progress_flag ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/guard.cc bitmask_type emergency_mutex emergency_buffer malloc dependents_used vptr thrown_size __cxa_allocate_dependent_exception __cxa_free_dependent_exception emergency_used dependents_buffer ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/eh_alloc.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=eh_alloc.lo get_new_handler _ZSt15get_new_handlerv ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/new_op.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=new_op.lo _ZNSt10bad_typeidD2Ev ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/bad_typeid.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=bad_typeid.lo _ZNSt10bad_typeidD0Ev ~bad_typeid _ZNKSt10bad_typeid4whatEv ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/guard_error.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=guard_error.lo _ZN9__gnu_cxx20recursive_init_errorD0Ev ~recursive_init_error _ZN9__gnu_cxx20recursive_init_errorD2Ev GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=pure.lo ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/pure.cc __cxa_pure_virtual __cxa_deleted_virtual contained_nonvirtual_p origin whole_object GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=dyncast.lo adjust_pointer<__cxxabiv1::(anonymous namespace)::vtable_prefix> ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/dyncast.cc whole_type whole_ptr vtable_prefix __cxa_bad_typeid __cxa_throw_bad_array_new_length ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/eh_aux_runtime.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=eh_aux_runtime.lo __cxa_throw_bad_array_length _ZN10__cxxabiv120__si_class_type_infoD2Ev _ZN10__cxxabiv120__si_class_type_infoD0Ev _ZN10__cxxabiv120__si_class_type_infoaSERKS0_ GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=si_class_type_info.lo _ZNK10__cxxabiv120__si_class_type_info11__do_upcastEPKNS_17__class_type_infoEPKvRNS1_15__upcast_resultE ~__si_class_type_info ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/si_class_type_info.cc _ZNK10__cxxabiv120__si_class_type_info12__do_dyncastElNS_17__class_type_info10__sub_kindEPKS1_PKvS4_S6_RNS1_16__dyncast_resultE _ZNK10__cxxabiv120__si_class_type_info20__do_find_public_srcElPKvPKNS_17__class_type_infoES2_ ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/eh_term_handler.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=eh_term_handler.lo __cxa_current_exception_type __cxa_demangle _ZN9__gnu_cxx27__verbose_terminate_handlerEv __builtin_fwrite fputs terminating __verbose_terminate_handler ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/vterminate.cc status GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=vterminate.lo __builtin_fputc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=eh_type.lo ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/eh_type.cc ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/eh_unex_handler.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=eh_unex_handler.lo ~bad_array_length GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=bad_array_length.lo _ZNSt16bad_array_lengthD0Ev _ZNSt16bad_array_lengthD2Ev ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/bad_array_length.cc _ZNKSt16bad_array_length4whatEv fake_num_cache_c _ZNSt6locale5_Impl13_S_id_collateE get_locale_mutex _M_init_facet<std::money_put<char> > fake_locale_Impl __mpcf facet_vec __mpct timepunct_cache_c _M_init_facet<std::time_get<char> > moneypunct_cf moneypunct_ct __facet name_vec _ZNSt6locale5_Impl11_S_id_ctypeE _M_init_facet<std::messages<char> > _ZNSt6locale5_Impl14_S_id_messagesE fake_num_put_c _M_init_facet<std::num_get<char> > fake_ctype_c fake_time_put_c ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/locale_init.cc fake_money_put_c _M_init_facet<std::numpunct<char> > fake_timepunct_c _M_init_facet<std::moneypunct<char, false> > __other_name _ZNSt6locale5_Impl10_S_id_timeE fake_time_cache_c GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=locale_init.lo fake_messages_c fake_num_get_c _ZNSt6locale5_Impl14_S_id_monetaryE _M_init_facet<std::codecvt<char, char, mbstate_t> > operator==<char, std::char_traits<char>, std::allocator<char> > _ZNSt6locale5_Impl19_S_facet_categoriesE fake_time_get_c _M_init_facet<std::time_put<char> > fake_money_get_c __npc fake_collate_c fake_locale _M_init_facet<std::ctype<char> > __tpc fake_codecvt_c _M_init_facet<std::money_get<char> > _ZNSt6locale5_ImplC2Em moneypunct_cache_cf fake_moneypunct_c _M_init_facet<std::num_put<char> > operator!=<char, std::char_traits<char>, std::allocator<char> > _M_init_facet<std::moneypunct<char, true> > _ZNSt6localeC2Ev c_locale_impl cache_vec _M_init_facet<std::__timepunct<char> > fake_money_cache_c name_c money_cache_cf numpunct_cache_c money_cache_ct _ZNSt6locale5_Impl13_S_id_numericE moneypunct_cache_ct _M_init_facet<std::collate<char> > fake_numpunct_c ~failure _ZNSt8ios_base7failureD2Ev ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/ios_failure.cc _ZNKSt8ios_base7failure4whatEv GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=ios_failure.lo _ZNSt8ios_base7failureD0Ev _M_msg _ZNSt8ios_base7failureC2ERKSs __table GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=ctype_configure_char.lo ctype_configure_char.cc __del _ZNSt5ctypeIcEC2EPKjbm _ZNSt5ctypeIcEC2EPiPKjbm collate_members.cc __cmp GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=collate_members.lo ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/globals_io.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=globals_io.lo fake_ostream fake_stdiobuf fake_filebuf fake_istream _ZNSdD0Ev GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=iostream-inst.lo _ZNSdD1Ev _ZSt7setfillIcESt8_SetfillIT_ES1_ ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/iostream-inst.cc _ZNSdD2Ev _ZNSdC2EPSt15basic_streambufIcSt11char_traitsIcEE _ZNSdC1Ev _ZNSdC1EPSt15basic_streambufIcSt11char_traitsIcEE setfill<char> _ZNSdC2Ev _ZNSt8numpunctIcED0Ev numeric_members.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=numeric_members.lo _ZNSt8numpunctIcED2Ev _ZNSirsEPFRSiS_E _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St12_Setiosflags _ZNSi3getERSt15basic_streambufIcSt11char_traitsIcEE _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE7_M_findIcEEN9__gnu_cxx11__enable_ifIXsrSt9__is_charIT_E7__valueEiE6__typeEPKS9_mS9_ _ZNSi3getEPclc _ZNSirsERb _ZNSirsERd _ZNSirsERe _ZNSirsERf _ZNSirsERi _ZNSirsERl _ZNSirsERm _ZNSirsERs _ZNSirsERt _ZNSirsERx _ZNSirsERy putback _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St8_SetfillIS3_E _ZSt2wsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_ _ZNSi4syncEv _ZNKSi6gcountEv _ZNSiC2EPSt15basic_streambufIcSt11char_traitsIcEE _M_extract<bool> _ZNSi10_M_extractIbEERSiRT_ _ZNSi10_M_extractIdEERSiRT_ _ZNSi10_M_extractIeEERSiRT_ _ZNSi10_M_extractIfEERSiRT_ _ZNSi10_M_extractIjEERSiRT_ _ZNSi10_M_extractIlEERSiRT_ _ZNSi10_M_extractImEERSiRT_ _ZNSi7getlineEPcl _ZNSi10_M_extractItEERSiRT_ _ZNSi10_M_extractIxEERSiRT_ _ZNSi10_M_extractIyEERSiRT_ _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St8_Setbase _ZNSi3getERc operator>><std::char_traits<char> > _M_extract<short unsigned int> _ZNSi4readEPcl _ZNSi6sentryC2ERSib _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_RS3_ ws<char, std::char_traits<char> > GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=istream-inst.lo _ZNSi5seekgESt4fposI9mbstate_tE _ZNSiC2Ev _ZNSi7putbackEc _ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Pa _ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Ph _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St14_Resetiosflags _ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Ra _ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Rh _ZNSi3getEPcl _ZNSi5ungetEv _M_extract<long double> _M_extract<long int> ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/istream-inst.cc _M_gcount _vptr.basic_istream __ng _M_extract<long long unsigned int> _ZNSi10_M_extractIPvEERSiRT_ _M_extract<void*> seekg tellg _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St13_Setprecision _ZNSi5seekgExSt12_Ios_Seekdir _ZNSiD0Ev __check_facet<std::num_get<char> > unget _ZNSirsEPFRSt9basic_iosIcSt11char_traitsIcEES3_E readsome _M_extract<long unsigned int> peek _ZNSi5tellgEv _ZNSiD1Ev _ZNSi3getEv _ZNSi3getERSt15basic_streambufIcSt11char_traitsIcEEc _ZNSirsERPv _ZNSirsEPSt15basic_streambufIcSt11char_traitsIcEE _M_extract<long long int> _ZNSi8readsomeEPcl _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St5_Setw __noskip _ZNSiD2Ev _ZNSirsERj _ZNSiC1Ev __this_sb _M_extract<double> _ZNSi4peekEv _M_extract<float> _ZNSiC1EPSt15basic_streambufIcSt11char_traitsIcEE _ZNSirsEPFRSt8ios_baseS0_E operator>> _M_extract<unsigned int> ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/ios_locale.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=ios_locale.lo xwrite st_blksize st_blocks _ZNSt14numeric_limitsIxE7epsilonEv __buffer _ZNSt12__basic_fileIcED2Ev dev_t nlink_t _ZNSt14numeric_limitsIxE10denorm_minEv fopen_mode errno st_uid _ZNSt12__basic_fileIcEC2EPi numeric_limits<long long int> _ZNSt14numeric_limitsIxE3minEv st_ctime st_nlink __c_mode st_gid ino_t __file st_size fstat st_mode _ZNSt14numeric_limitsIxE13signaling_NaNEv blkcnt_t FsVirtID mode_t st_atime lseek st_dev basic_file.cc fdopen st_mtime _ZNSt14numeric_limitsIxE8infinityEv _ZNSt14numeric_limitsIxE3maxEv _ZNSt14numeric_limitsIxE9quiet_NaNEv uid_t blksize_t _ZNSt14numeric_limitsIxE11round_errorEv st_ino gid_t GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=basic_file.lo GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=messages_members.lo messages_members.cc _ZNSt12out_of_rangeD0Ev _ZNSt13runtime_errorC2ERKSs _ZNSt11logic_errorD0Ev _ZNSt12domain_errorC2ERKSs _ZNSt16invalid_argumentD2Ev _ZNSt12out_of_rangeD2Ev ~domain_error ../../../../../gcc-4.9.1/libstdc++-v3/src/c++98/stdexcept.cc _ZNSt15underflow_errorC2ERKSs _ZNSt11range_errorD0Ev _ZNKSt11logic_error4whatEv ~runtime_error _ZNSt12length_errorD0Ev _ZNSt12length_errorD2Ev _ZNSt14overflow_errorC2ERKSs _ZNSt12domain_errorD2Ev ~range_error ~length_error _ZNSt11logic_errorD2Ev _ZNSt15underflow_errorD0Ev _ZNSt11logic_errorC2ERKSs _ZNSt12length_errorC2ERKSs _ZNSt13runtime_errorD0Ev _ZNSt14overflow_errorD0Ev ~logic_error GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=stdexcept.lo _ZNSt16invalid_argumentD0Ev _ZNSt11range_errorD2Ev ~out_of_range ~invalid_argument _ZNSt13runtime_errorD2Ev ~overflow_error _ZNSt16invalid_argumentC2ERKSs _ZNSt15underflow_errorD2Ev _ZNSt11range_errorC2ERKSs _ZNKSt13runtime_error4whatEv _ZNSt12out_of_rangeC2ERKSs ~underflow_error _ZNSt12domain_errorD0Ev _ZNSt14overflow_errorD2Ev _ZNSt14numeric_limitsIdE11round_errorEv c++locale.cc numeric_limits<double> _ZNSt14numeric_limitsIdE3maxEv _ZNSt14numeric_limitsIeE3maxEv __overflow _ZNSt14numeric_limitsIfE7epsilonEv numeric_limits<float> _ZNSt14numeric_limitsIfE3maxEv _ZNSt14numeric_limitsIeE3minEv category_names _ZNSt6locale13_S_categoriesE __sanity sscanf _ZNSt14numeric_limitsIdE8infinityEv _ZNSt14numeric_limitsIfE8infinityEv _ZNSt14numeric_limitsIdE13signaling_NaNEv _ZNSt14numeric_limitsIeE13signaling_NaNEv numeric_limits<long double> _ZNSt14numeric_limitsIfE13signaling_NaNEv _ZNSt14numeric_limitsIdE10denorm_minEv _ZNSt14numeric_limitsIeE8infinityEv _ZNSt14numeric_limitsIdE9quiet_NaNEv _ZNSt14numeric_limitsIfE10denorm_minEv strtof _ZNSt14numeric_limitsIeE10denorm_minEv _ZNSt14numeric_limitsIfE9quiet_NaNEv _ZNSt14numeric_limitsIeE7epsilonEv _ZNSt14numeric_limitsIeE9quiet_NaNEv _ZNSt14numeric_limitsIfE11round_errorEv _ZNSt14numeric_limitsIeE11round_errorEv _ZNSt14numeric_limitsIdE3minEv _ZNSt14numeric_limitsIdE7epsilonEv _ZNSt14numeric_limitsIfE3minEv GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=c++locale.lo GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=time_members.lo __llen time_members.cc GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=functional.lo ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11/functional.cc ~bad_function_call _ZNSt17bad_function_callD2Ev _ZNKSt17bad_function_call4whatEv _ZNSt17bad_function_callD0Ev GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=snprintf_lite.lo __errlen __throw_insufficient_space __val2 ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11/snprintf_lite.cc __concat_size_t __bufsize _ZN9__gnu_cxx15__concat_size_tEPcmm _ZN9__gnu_cxx26__throw_insufficient_spaceEPKcS1_ memory_order_acquire memory_order_acq_rel _ZNSt12future_errorD0Ev __cxa_atexit memory_order_consume memory_order_seq_cst GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=future.lo __future_category_instance _ZNKSt12future_error4codeEv ~future_error_category memory_order_relaxed ~future_error __fec _ZNSt12future_errorD2Ev ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11/future.cc _ZNKSt12future_error4whatEv __dso_handle memory_order_release memory_order __cond ~system_error_category ~generic_error_category _ZNKSt14error_categoryneERKS_ _ZNKSt14error_category23default_error_conditionEi ~system_error operator< ../../../../../gcc-4.9.1/libstdc++-v3/src/c++11/system_error.cc _ZNKSt14error_category10equivalentERKSt10error_codei _ZNKSt14error_category7messageEi _ZNKSt12system_error4codeEv generic_category_instance _vptr.error_category _ZNKSt14error_category10equivalentEiRKSt15error_condition _ZNKSt14error_categoryltERKS_ _ZNKSt14error_category4nameEv _ZNSt12system_errorD0Ev _ZNKSt14error_categoryeqERKS_ system_category ~error_category _GLOBAL__sub_I__ZNSt14error_categoryD2Ev system_category_instance equivalent __code _ZNSt12system_errorD2Ev _ZNSt14error_categoryD0Ev _ZSt15system_categoryv _ZNSt14error_categoryaSERKS_ GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=system_error.lo _ZSt15set_new_handlerPFvvE ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/new_handler.cc set_new_handler __new_handler prev_handler GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=new_handler.lo GNU C++ 4.9.1 -mtune=generic -march=pentiumpro -g -O2 -std=gnu++11 -fno-implicit-templates -ffunction-sections -fdata-sections -frandom-seed=bad_array_new.lo _ZNKSt20bad_array_new_length4whatEv ../../../../gcc-4.9.1/libstdc++-v3/libsupc++/bad_array_new.cc _ZNSt20bad_array_new_lengthD0Ev ~bad_array_new_length _ZNSt20bad_array_new_lengthD2Ev DEMANGLE_COMPONENT_OPERATOR D_PRINT_DEFAULT DEMANGLE_COMPONENT_TYPEINFO_NAME d_template_arg DEMANGLE_COMPONENT_DEFAULT_ARG d_make_comp d_builtin_type_print hold_current d_make_extended_operator d_bare_function_type d_make_character d_cv_qualifiers DEMANGLE_COMPONENT_RVALUE_REFERENCE D_PRINT_INT full_expansion d_print_callback DEMANGLE_COMPONENT_CONST d_local_name estimate pstart simple d_identifier d_print_mod_list d_init_info is_expression d_compact_number next_sub d_make_ctor gnu_v3_base_object_ctor GNU C 4.9.1 -mtune=generic -march=pentiumpro -g -O2 s_builtin DEMANGLE_COMPONENT_RESTRICT_THIS d_class_enum_type DEMANGLE_COMPONENT_VTABLE d_print_cast DEMANGLE_COMPONENT_UNARY current_template d_growable_string demangle_component_type is_ctor_dtor_or_conversion comb_type DEMANGLE_COMPONENT_BINARY d_lambda DEMANGLE_COMPONENT_DECLTYPE DEMANGLE_COMPONENT_THUNK DEMANGLE_COMPONENT_BINARY_ARGS s_name op_is_new_cast DEMANGLE_COMPONENT_NULLARY d_info member_fn d_pointer_to_member_type did_subs template_decl demangled DEMANGLE_COMPONENT_REFERENCE_THIS next_saved_scope derived_type d_ctor_dtor_name D_PRINT_FLOAT d_add_substitution is_conversion DEMANGLE_COMPONENT_VECTOR_TYPE DEMANGLE_COMPONENT_ARRAY_TYPE d_java_resource discrim DEMANGLE_COMPONENT_SUB_STD DCT_GLOBAL_DTORS DEMANGLE_COMPONENT_TAGGED_NAME realloc d_print_info gnu_v3_complete_object_ctor DEMANGLE_COMPONENT_TYPEINFO d_last_char simple_expansion DEMANGLE_COMPONENT_FUNCTION_TYPE DEMANGLE_COMPONENT_GLOBAL_DESTRUCTORS d_print_saw_error d_template_param num_subs d_operator_name DEMANGLE_COMPONENT_TEMPLATE_ARGLIST d_print_expr_op DEMANGLE_COMPONENT_CTOR d_fill_extended_operator DEMANGLE_COMPONENT_VTT java_name d_expression_1 d_append_buffer peek_next newalc DCT_GLOBAL_CTORS d_standard_sub_info DEMANGLE_COMPONENT_UNNAMED_TYPE d_make_operator need d_print_init d_demangle_callback standard_subs DEMANGLE_COMPONENT_CHARACTER gnu_v3_unified_dtor DEMANGLE_COMPONENT_IMAGINARY DEMANGLE_COMPONENT_QUAL_NAME d_expr_primary cplus_demangle_builtin_types d_backtrack flush_count DEMANGLE_COMPONENT_VOLATILE_THIS hold_dpm DEMANGLE_COMPONENT_TLS_WRAPPER accum hold_dpt d_make_demangle_mangled_name DEMANGLE_COMPONENT_HIDDEN_ALIAS d_unnamed_type DEMANGLE_COMPONENT_TEMPLATE DEMANGLE_COMPONENT_COVARIANT_THUNK gnu_v3_deleting_dtor d_template_args D_PRINT_LONG_LONG need_space terminator D_PRINT_UNSIGNED_LONG_LONG full_len DEMANGLE_COMPONENT_ARGLIST d_call_offset d_growable_string_resize d_growable_string_append_buffer num_scopes DEMANGLE_COMPONENT_LITERAL DEMANGLE_COMPONENT_FIXED_TYPE DEMANGLE_COMPONENT_COMPOUND_NAME d_print_flush d_fill_dtor d_append_num send java_len s_ctor verbose hold_last_name printed DEMANGLE_COMPONENT_REFTEMP DEMANGLE_COMPONENT_CONST_THIS second DEMANGLE_COMPONENT_TYPEINFO_FN s_unary_num d_make_default_arg pdpm d_append_string d_print_java_identifier saved_templates d_get_saved_scope gnu_v3_dtor_kinds d_prefix D_PRINT_BUFFER_LENGTH d_count_templates_scopes DCT_MANGLED d_expression d_unqualified_name mod_inner DEMANGLE_COMPONENT_CLONE d_info_checkpoint DCT_TYPE simple_len third d_array_type next_copy_template DEMANGLE_COMPONENT_COMPLEX DEMANGLE_COMPONENT_VOLATILE d_make_template_param DEMANGLE_COMPONENT_PACK_EXPANSION d_make_dtor s_string DEMANGLE_COMPONENT_JAVA_RESOURCE gnu_v3_base_object_dtor d_save_scope DEMANGLE_COMPONENT_CAST d_clone_suffix demangle_builtin_type_info num_templates DEMANGLE_COMPONENT_TRANSACTION_CLONE d_fill_name d_number s_operator temps d_saved_scope top_level d_abi_tags opaque d_print_comp d_make_sub d_print_template can_subst d_make_builtin_type d_parmlist D_PRINT_VOID DEMANGLE_COMPONENT_BUILTIN_TYPE DEMANGLE_COMPONENT_TEMPLATE_PARAM s_character demangle_operator_info gnu_v3_object_dtor_group d_index_template_argument set_last_name d_vector_type d_ref_qualifier DEMANGLE_COMPONENT_VIRTUAL_THUNK gnu_v3_ctor_kinds DEMANGLE_COMPONENT_LAMBDA d_nested_name has_return_type s_binary peek2 recurse_left_right demangle_callbackref d_growable_string_init demangle_component d_make_function_param d_checkpoint s_fixed d_special_name DEMANGLE_COMPONENT_RVALUE_REFERENCE_THIS was_expression D_PRINT_UNSIGNED d_make_name num_copy_templates gnu_v3_complete_object_dtor next_comp DEMANGLE_COMPONENT_TRINARY d_print_function_type DEMANGLE_COMPONENT_VENDOR_TYPE_QUAL d_make_empty palc d_append_char DEMANGLE_COMPONENT_TYPED_NAME D_PRINT_BOOL d_print_array_type num_saved_scopes DEMANGLE_COMPONENT_POINTER modifier DEMANGLE_COMPONENT_LOCAL_NAME pack_index D_PRINT_LONG cplus_demangle_operators DEMANGLE_COMPONENT_NONTRANSACTION_CLONE need_paren new_id DEMANGLE_COMPONENT_REFERENCE DEMANGLE_COMPONENT_TRINARY_ARG1 DEMANGLE_COMPONENT_TRINARY_ARG2 DEMANGLE_COMPONENT_DTOR DEMANGLE_COMPONENT_GUARD DEMANGLE_COMPONENT_VENDOR_TYPE newbuf s_number mods hold_modifiers DEMANGLE_COMPONENT_FUNCTION_PARAM d_print_subexpr d_source_name d_demangle set_last_name_len d_find_pack DEMANGLE_COMPONENT_TLS_INIT s_extended_operator gnu_v3_unified_ctor gnu_v3_object_ctor_group DEMANGLE_COMPONENT_GLOBAL_CONSTRUCTORS d_growable_string_callback_adapter d_discriminator DEMANGLE_COMPONENT_NUMBER demangle_failure __gcclibcxx_demangle_callback container d_exprlist DEMANGLE_COMPONENT_INITIALIZER_LIST d_print_error d_pack_length cp-demangle.c adpm output_buffer DEMANGLE_COMPONENT_RESTRICT d_print_mod d_number_component d_function_type options DEMANGLE_COMPONENT_EXTENDED_OPERATOR rqual gnu_v3_complete_object_allocating_ctor need_template_restore typed_name DEMANGLE_COMPONENT_LITERAL_NEG DEMANGLE_COMPONENT_NAME DEMANGLE_COMPONENT_CONSTRUCTION_VTABLE DEMANGLE_COMPONENT_JAVA_CLASS d_mangled_name d_fill_ctor DEMANGLE_COMPONENT_PTRMEM_TYPE num_comps D_PRINT_UNSIGNED_LONG allocation_failure d_lookup_template_argument was_conversion s_dtor operand complex double USItype DWunion complex float DWstruct /opt/MeetiXOSProject/temp/build-gcc/i686-mx/libgcc complex long double __udivdi3 ../../../gcc-4.9.1/libgcc/libgcc2.c __udivmoddi4 GNU C 4.9.1 -mtune=generic -march=pentiumpro -g -g -g -O2 -O2 -O2 -fbuilding-libgcc -fno-stack-protector -fpic -fexceptions -fnon-call-exceptions -fvisibility=hidden UDItype __umoddi3 DW_OP_GNU_addr_index lsda_encoding DW_OP_HP_unknown X86_TUNE_MEMORY_MISMATCH_STALL DW_OP_lit15 DW_CFA_lo_user DW_OP_lit17 X86_TUNE_READ_MODIFY DW_OP_HP_unmod_range X86_TUNE_ALWAYS_FANCY_MATH_387 DW_OP_breg4 uword X86_TUNE_SSE_PACKED_SINGLE_INSN_OPTIMAL DW_OP_GNU_encoded_addr X86_TUNE_ZERO_EXTEND_WITH_AND uw_install_context_1 X86_TUNE_USE_BT DW_OP_GNU_regval_type DW_OP_lit0 DW_OP_lit1 DW_OP_lit2 DW_OP_lit3 DW_OP_lit4 DW_OP_lit5 DW_OP_lit6 DW_OP_lit8 DW_OP_lit9 old_rs DW_OP_call_ref DW_OP_GNU_const_index X86_TUNE_USE_HIMODE_FIOP X86_TUNE_PARTIAL_FLAG_REG_STALL X86_TUNE_PUSH_MEMORY X86_TUNE_INTER_UNIT_MOVES_TO_VEC _Unwind_GetPtr X86_TUNE_MOVE_M1_VIA_OR REG_SAVED_VAL_OFFSET DW_CFA_def_cfa DW_CFA_MIPS_advance_loc8 X86_TUNE_AVOID_LEA_FOR_ADDR X86_TUNE_AVX256_UNALIGNED_STORE_OPTIMAL DW_CFA_set_loc execute_stack_op unused_rs cfa_exp DW_CFA_offset DW_OP_abs new_rs DW_OP_reg11 DW_OP_reg12 DW_OP_reg13 DW_OP_reg14 DW_OP_reg15 DW_OP_reg17 DW_OP_reg18 DW_OP_drop outer_cfa DW_CFA_register DW_OP_HP_tls DW_CFA_val_offset X86_TUNE_PROMOTE_QI_REGS X86_TUNE_USE_SIMODE_FIOP X86_TUNE_MOVX signal_frame X86_TUNE_SPLIT_MEM_OPND_FOR_FP_CONVERTS DW_OP_reg20 DW_OP_reg21 DW_OP_reg22 DW_OP_reg23 DW_OP_mul DW_OP_reg25 DW_OP_reg26 DW_OP_reg27 DW_OP_reg29 extract_cie_info DW_OP_nop DW_OP_not dwarf_location_atom DW_OP_GNU_implicit_pointer DW_OP_plus DW_OP_const2s DW_OP_xor DW_CFA_def_cfa_offset DW_OP_piece DW_OP_reg30 DW_OP_reg31 dwarf_fde stop_code X86_TUNE_VECTORIZE_DOUBLE eh_ptr X86_TUNE_SOFTWARE_PREFETCHING_BENEFICIAL saved X86_TUNE_AVOID_VECTOR_DECODE ../../../gcc-4.9.1/libgcc/unwind-dw2.c _Unwind_Personality_Fn DW_CFA_val_offset_sf saw_z X86_TUNE_SHIFT1 uw_update_context_1 X86_TUNE_SSE_SPLIT_REGS DW_OP_deref stack_elt X86_TUNE_INTER_UNIT_CONVERSIONS DW_OP_GNU_deref_type read_2s X86_ARCH_CMPXCHG8B ix86_tune_indices X86_TUNE_SSE_PARTIAL_REG_DEPENDENCY CFA_EXP DW_OP_const2u dwarf_cie cur_context DW_CFA_def_cfa_offset_sf DW_OP_breg0 X86_TUNE_REASSOC_INT_TO_PARALLEL X86_TUNE_FUSE_CMP_AND_BRANCH_64 DW_OP_breg3 X86_TUNE_DOUBLE_PUSH X86_TUNE_FUSE_ALU_AND_BRANCH DW_OP_HP_mod_range _Unwind_GetGRPtr X86_TUNE_INTEGER_DFMODE_MOVES X86_ARCH_BSWAP REG_SAVED_OFFSET pc_begin X86_TUNE_SSE_UNALIGNED_STORE_OPTIMAL target_cfa DW_OP_PGI_omp_thread_num _Unwind_Trace_Fn X86_TUNE_DOUBLE_POP X86_TUNE_USE_FFREEP uw_update_context DW_OP_consts DW_OP_stack_value DW_OP_constu uw_identify_context DW_OP_GNU_entry_value DW_OP_form_tls_address DW_OP_plus_uconst match_handler X86_TUNE_UNROLL_STRLEN sword DW_OP_shra DW_OP_const4s _Unwind_ForcedUnwind DW_OP_dup X86_TUNE_LCP_STALL REG_SAVED_REG DW_OP_eq REG_SAVED_EXP frame_state_reg_info _Unwind_Find_FDE DW_OP_xderef_size DW_OP_call2 _Unwind_GetGR CFA_REG_OFFSET X86_TUNE_PAD_SHORT_FUNCTION DW_OP_call_frame_cfa DW_CFA_advance_loc X86_TUNE_SSE_UNALIGNED_LOAD_OPTIMAL tmp_sp op_ptr X86_TUNE_PROLOGUE_USING_MOVE DW_OP_ge DW_OP_lit20 REG_SAVED_VAL_EXP DW_OP_lit24 DW_OP_HP_fltconst4 cfa_how DW_OP_fbreg DW_OP_HP_fltconst8 DW_OP_gt X86_TUNE_USE_SAHF X86_TUNE_AVOID_MEM_OPND_FOR_CMOVE X86_TUNE_ADJUST_UNROLL CFA_UNSET uw_advance_context _Unwind_GetIP execute_cfa_program no_push DW_OP_reg7 DW_OP_breg14 X86_TUNE_USE_LEAVE DW_OP_breg15 X86_TUNE_USE_INCDEC X86_ARCH_XADD X86_TUNE_SSE_LOAD0_BY_PXOR DW_CFA_hi_user DW_OP_const8s DW_OP_const8u stmp X86_TUNE_SLOW_IMUL_IMM8 DW_CFA_expression utmp DW_OP_GNU_parameter_ref X86_TUNE_SCHEDULE X86_TUNE_USE_XCHGB DW_OP_and ubyte this_context DW_OP_breg22 DW_CFA_restore X86_TUNE_EPILOGUE_USING_MOVE X86_TUNE_FAST_PREFIX op_end state_in cfa_reg X86_TUNE_FUSE_CMP_AND_BRANCH_SOFLAGS outer_ra DW_OP_lo_user _Unwind_IsExtendedContext X86_TUNE_GENERAL_REGS_SSE_SPILL DW_OP_pick DW_OP_breg1 DW_OP_breg2 X86_TUNE_DOUBLE_WITH_ADD DW_OP_breg5 DW_OP_breg6 DW_OP_breg7 DW_OP_breg8 DW_OP_breg9 stop read_1s read_1u DW_OP_HP_is_value X86_TUNE_READ_MODIFY_WRITE _Unwind_SetSpColumn retaddr_column _Unwind_Stop_Fn _Unwind_Backtrace DW_CFA_same_value X86_TUNE_NOT_VECTORMODE _Unwind_SetGRPtr DW_OP_bregx DW_OP_le reg_or_offset read_2u DW_OP_lt _Unwind_FrameState augmentation DW_CFA_restore_extended DW_OP_minus CIE_delta DW_OP_implicit_value _Unwind_FindEnclosingFunction X86_TUNE_SINGLE_POP DW_CFA_def_cfa_expression uw_init_context_1 DW_OP_GNU_uninit DW_CFA_restore_state X86_TUNE_NOT_UNPAIRABLE X86_TUNE_QIMODE_MATH X86_TUNE_USE_VECTOR_CONVERTS X86_TUNE_SINGLE_PUSH X86_TUNE_PARTIAL_REG_STALL DW_OP_lit30 DW_OP_ne read_4s read_4u X86_ARCH_CMOV DW_OP_GNU_convert _Unwind_DebugHook DW_OP_xderef DW_OP_skip DW_OP_GNU_reinterpret DW_OP_const1s DW_OP_const1u init_dwarf_reg_size_table X86_TUNE_USE_MOV0 X86_TUNE_SSE_TYPELESS_STORES DW_OP_or read_pointer REG_UNSAVED _Unwind_ForcedUnwind_Phase2 X86_TUNE_USE_VECTOR_FP_CONVERTS DW_OP_lit10 DW_OP_lit11 DW_OP_lit12 DW_OP_lit13 DW_OP_lit14 X86_TUNE_PARTIAL_REG_DEPENDENCY DW_OP_lit16 DW_OP_lit18 DW_OP_lit19 _Unwind_SetSignalFrame DW_CFA_advance_loc1 DW_CFA_advance_loc2 DW_CFA_advance_loc4 uw_frame_state_for X86_TUNE_LAST DW_CFA_GNU_negative_offset_extended DW_OP_breg10 DW_OP_breg11 DW_OP_breg12 DW_OP_breg13 DW_OP_breg16 DW_OP_breg17 DW_OP_breg18 DW_OP_breg19 DW_OP_lit21 DW_OP_lit22 DW_OP_lit23 X86_TUNE_SLOW_IMUL_IMM32_MEM DW_OP_lit25 DW_OP_lit26 DW_OP_lit27 DW_OP_lit28 DW_OP_lit29 DW_OP_GNU_const_type __frame_state_for DW_CFA_undefined pc_target _Unwind_RaiseException_Phase2 DW_OP_mod DW_OP_breg20 DW_OP_breg21 regs DW_OP_breg23 DW_OP_breg24 DW_OP_breg25 DW_OP_breg26 DW_OP_breg27 DW_OP_breg28 DW_OP_breg29 DW_OP_lit31 insn_ptr X86_TUNE_AVX256_UNALIGNED_LOAD_OPTIMAL by_value X86_TUNE_ACCUMULATE_OUTGOING_ARGS DW_CFA_def_cfa_register read_8s read_8u orig_context _Unwind_IsSignalFrame DW_OP_breg30 DW_OP_breg31 _Unwind_SetGRValue frame_state DW_OP_push_object_address X86_TUNE_BRANCH_PREDICTION_HINTS DW_OP_over X86_TUNE_AVX128_OPTIMAL DW_CFA_offset_extended_sf DW_OP_swap DW_CFA_remember_state DW_OP_reg10 DW_OP_reg16 DW_OP_reg19 DW_CFA_GNU_window_save DW_OP_neg DW_CFA_offset_extended DW_OP_bra X86_TUNE_OPT_AGU _Unwind_Get_Unwind_Context_Reg_Val X86_TUNE_HIMODE_MATH DW_OP_reg0 DW_OP_reg1 DW_OP_reg2 DW_OP_reg3 DW_OP_reg4 DW_OP_reg5 DW_OP_reg6 personality DW_OP_reg8 DW_OP_reg9 DW_OP_GNU_push_tls_address get_cie DW_OP_const4u X86_TUNE_SPLIT_LONG_MOVES DW_CFA_val_expression DW_OP_call4 X86_TUNE_PROMOTE_HIMODE_IMUL X86_TUNE_EXT_80387_CONSTANTS _Unwind_SpTmp DW_OP_regx X86_TUNE_SINGLE_STRINGOP sp_slot DW_OP_reg24 X86_TUNE_FOUR_JUMP_LIMIT DW_OP_reg28 CIE_id GNU C 4.9.1 -mtune=generic -march=pentiumpro -g -g -g -O2 -O2 -O2 -fbuilding-libgcc -fno-stack-protector -fpic -fexceptions -fvisibility=hidden X86_TUNE_REASSOC_FP_TO_PARALLEL trace_argument data_align X86_TUNE_MISALIGNED_MOVE_STRING_PRO_EPILOGUES initial X86_ARCH_LAST next_fde ix86_arch_indices _Unwind_GetCFA X86_TUNE_PAD_RETURNS X86_TUNE_PROMOTE_HI_REGS DW_OP_bit_piece REG_UNDEFINED DW_OP_shl DW_OP_deref_size DW_OP_shr code_align DW_CFA_GNU_args_size X86_TUNE_FUSE_CMP_AND_BRANCH_32 dwarf_eh_bases dbase X86_TUNE_INTER_UNIT_MOVES_FROM_VEC X86_TUNE_USE_CLTD DW_OP_div X86_TUNE_PROMOTE_QIMODE DW_CFA_nop _Unwind_Get_Unwind_Word DW_OP_rot _Unwind_GRByValue dwarf_call_frame_info presult insn_end stop_argument DW_CFA_def_cfa_sf X86_ARCH_CMPXCHG DW_OP_addr DW_OP_hi_user DW_OP_lit7 binary_search_unencoded_fdes fde_insert erratic pc_array y_encoding this_cie unseen_objects fde_mixed_encoding_compare __gthread_mutex_lock __register_frame_table probe linear ../../../gcc-4.9.1/libgcc/unwind-dw2-fde.c fde_accumulator last_cie cur_count __deregister_frame_info_bases __register_frame_info end_fde_sort uaddr get_cie_encoding fini fde_compare accu start_fde_sort from_array __gthread_mutex_unlock __register_frame_info_table_bases unhandled_fdes pc_range binary_search_single_encoding_fdes frame_heapsort fde_vector fde_unencoded_compare y_ptr binary_search_mixed_encoding_fdes object_mutex marker __register_frame_info_bases frame_downheap chain_end base_from_object fde_compare_t __register_frame linear_search_fdes fde_merge fde2 fde_split classify_object_over_fdes init_object search_object last_fde mixed_encoding x_encoding add_fdes __deregister_frame_info __register_frame_info_table fde_single_encoding_compare orig_data sorted this_fde x_ptr __deregister_frame get_fde_encoding �� P�0� P        ��� R��/� W/�0� �R�        ��� 0���� Q�� qy��0� Q        �� R�,� p        ��� 0���.� V.�/� w /�0� �R        0�>� P>�y� Vy�{� �P�        0�G� RG�x� Sx�{� �R�        0�G� QG�z� Wz�{� �Q�        ���� P��e� �P�e�w� Pw��� �P�        ���� R��ߑ �Lߑ� R�� �L�� R��� �L��� R�� �L�"� R"�N� �LN�S� RS�[� �L[�d� Rd�e� �Le�|� R|��� �L        ���� Q��ۑ Sۑߑ Pߑ� Q�� S��� Q���� S��
� Q
�� V�� P�&� Q&�N� VN�V� QV�[� S[�d� Qd�e� Ve�� Q��� S���� P        ���� Q��ő Vőߑ �Q�ߑ
� Q
�� V�&� Q&�N� VN�d� Qd�e� Ve��� Q        ��ߑ R�� R��� R�� RS�[� R|��� R        0�N� S        0�A� QA�C� qy�C�N� Q        7�I� RI�N� s        0�N� U        e�z� Qz��� V���� p|�        ��ƒ Pƒْ �P�ْ�� P���� �P���� P        ���� R���� �R�ْ� R��� �R���� R�� �R��� R�� �R�        ��ʒ Sʒϒ Pْ� S         �8� P8��� W���� �P����� W���� �P�         �8� R8��� U���� �R����� U���� �R�         �8� Q8�v� �\v�|� q |��� �\        8�D� V        r�|� P        g�q� R���� R        8��� V���� V        8�D� 0�D�a� Qa�c� qy�c�q� Q���� Q        W�m� Pm�q� v���� P���� v        8�D� 0�D�q� R���� R        ���� P��� �P�        ��ē Rē̓ �R�̓� R�� �R���� R�� � �R� �� R�� �R�        �� P�j� Wj��� �P���� W�� �P�        �-� R-�8� U8�p� Vp��� R���� R���� P��� V�� R        �-� Q-�� �\        ���� W�� W        >�L� RL�R� vR�j� U��� R        G�V� s�V�^� R^�d� t d�j� s�        G�j� V        G�L� RL�R� vR�j� U        G�j� W        ���� R        ���� Q���� qy����� Q        ���� S        ���� W        ���� ��           ���� P        ��� Q�� qy���� Q        ה�� S        ��� W        ���� 3�N�p� P���� 1���ŗ Pҗ�� P%�/� 0�k�u� 3�        ���� P���� �@��� ��=�S� PS�[� R[��� ������ pp��� ��        ��R� 0���� 0�/�Q� 0�Q�_� P_��� R��,� W,�/� v p "�/�u� Wu�}� 0�Й� W�� R        ^�c� Pc�Ė S�� S���� W��Ř PŘg� VЙ�� V        ���� V��N� 0����� 0���� 0�/�?� 0�?�I� PI��� V��u� ��u�}� P}��� VЙ� ��        ���� P��I� V��� V/�?� V        ���� S��R� 0����� S��� 0�%�k� 0�k�u� Su��� 0�Й� 0�        z��� ���� ��        `�f� Q�S�        ���� �   ���� �           ���� �   ���� �           ���� ��   ���� ��           ���� ����� P        7�G� U��� U/��� Uu��� U        ��G� W��� W/��� W��u� ���u��� WЙ� ���        ��Ė S        ���� �]��Ɩ U        ��G� 0���� 0�/��� 0�Й� 0�        Ɩݖ �@�ݖ�� P��� t �G� �@���� �@�/��� �@����� R���� �@�Й� �@�        Ɩ͖ P͖� U        Ɩі �]і� S        ƖG� 0���� 0�/��� 0�Й� 0�        �� �D��� P�� t �G� �D���� �D�/��� �D���Ř RŘ�� �D�Й� �D�        �� P�� U�� Q        ��� �]��� S        �G� 0���� 0�/��� 0�Й� 0�         �G� S��� S/��� Su��� S         �1� Q1�3� qy�3�G� Q��� Q/��� Qu��� Q        '�G� R��� R/�Q� RQ��� su�}� R}��� s         �G� U��� U/��� Uu��� U        D�\� P        ��u� ��Й� ��        [��� 0���9� ��;�g� ��Й� ��        [�g� 0�Й�� 0�        ��� �        �� �H�        �� R�� �@        ���� R���	 �@ �T"�        �� U        ��� ��            ��� R        ���� 0���� Q�� qy��� Q        �� S        ���� 0���� U        v��� �        v��� ��        v��� ��        v��� �        ,�g� Sg��� u��� u        >�A� PA�H� spH�� uD        [�]� P        ]�s� P        ]�s� p0�        Κ� P        6�M� �         6�E� PE�V� �        }��� P        �� P,�6� P        �� R�'� sP�,�6� R        �� r0,�6� r0        U�x� s         ���� � ���� p|�        ���� � #����� P        ؜�� S���� �         �� P��� s����� � #�        �,� �         �0� �        L�O� s�O��� V���� u#����� t#���Ɲ V        a�j� P���� P        V��� V���� ����� V���� �        V�{� ����� �        V�`� P        h�{� �        h��� V���� �        h�m� Sm�t� �         m��� 1�        m�� S��� �         m�t� st�w� P        ��О 0�О� 1��f� 0�        ���� P        ڞ� 1�        ڞ� R        ڞ� r        �� 1�:�C� 1�H�V� 1�        �� S:�<� S>�C� S        �� s�:�<� s�>�C� s�        �� s        )�:� 1�C�H� 1�V�f� 1�        )�7� QC�G� Q        )�7� q�C�G� q�        )�-� q        ~��� S���� u���� t��� S�� u�� t�4� S4�6� u6�@� S@�N� uN�P� SP�^� u        ��ǟ P        ��� 1�2�;� 1�@�N� 1�        ��� V2�;� V@�N� V        ��� v�2�;� v�@�N� v�        ��� v        �2� 1�;�@� 1�N�^� 1�        �2� V;�@� VN�^� V        �2� v�;�@� v�N�^� v�        �"� v        `�y� 0���Š 0�Š� 4��Y� 0�        ���� P���� t ���� t        Ϡ� 4�        Ϡ۠ R        Ϡ֠ r        ��� 1�-�6� 1�;�I� 1�        ��� S-�/� S1�6� S        ��� s�-�/� s�1�6� s�        ���� s        �-� 1�6�;� 1�I�Y� 1�        �'� Q6�:� Q        �'� q�6�:� q�        �� q        `�� 0����� 0���ѡ 4�ѡI� 0�        ���� P        ��ѡ 4�        ��ˡ R        ��ơ r        ��� 1��&� 1�+�9� 1�        ��� S�� S!�&� S        ��� s��� s�!�&� s�        �� s        	�� 1�&�+� 1�9�I� 1�        	�� W&�+� W9�I� W        	�� w�&�+� w�9�I� w�        	�� w        P�p� �         P�l� �        ���� s���� V�� u#��� t#��� V        ]�c� R        ���� P        ˣף P        ˣң p        �9� 0����� 0�ɤФ 0��D� 0�        �!� v v <"#x        �9� Sɤˤ SˤФ u�/� S/�1� u1�=� S=�D� u        ˤФ 1���� 1�-�6� 1�        ˤФ V��� V-�6� V        ˤФ v���� v�-�6� v�        ���� v        �-� 4�6�D� 4�        �'� Q6�:� Q        �'� q�6�:� q�        �� q        C�L� Q        C�G� q        P��� u`����� t\���Ĥ u`�ĤŤ t\�        p�x� P        ��Ť 1�        ���� P        ���� p        r��� 0���� 0�:�<� 0�@�j� 0�{��� 0�        {��� W��
� W
�� Q��� W        {��� P��� P        �� P        ���� 1�        ��
� W
�� Q��� W        ��� P        %�:� 1�        %�1� R        %�,� r        V�j� 1�{��� 1�        V�e� V{�}� V��� V        V�e� v�{�}� v���� v�        V�Z� v        ���� Q���� Q        ���� q����� q�        ���� q        ��ť u`�ťƥ t\�ƥ�� u`����� t\�        ���� P        ۥ�� 1�        ۥ� P        ۥ� p        �� S��ӧ Sӧէ uէڧ Sڧ� u�� S��� u���� S��� u        �� u���� u���� u        �� V���� V��ѧ V�� V        ��� P        �� S��ӧ Sӧէ uէڧ Sڧ� u�� S��� u���� S��� u        �� u���� u���� u        ��� P        ��� u        ��� S        ��� V        	�� 1�        	�� R        	�� r        ���� 1�ѧߧ 1�        ���� Vѧߧ V        ���� v�ѧߧ v�        ���� v        ��ѧ 1��� 1�        ��˧ Q���� Q        ��˧ q����� q�        ���� q        �S� u`�S�T� t\�T��� u`����� t\�        9�A� P        k��� 1�        k�w� P        k�r� p        )�@�
 v v <"�X�h� v p "����� v p "�        2�R� SX��� S        6��� :�        6�R� SX��� S        X��� :�        X��� S        J�W� P        Ш� � �� S�� � �J� S        Ш� ��� P�� ��� P�J� �        ި� V�� V�J� V        �� v� �� v�         �� V�J� V        �� W�J� W        �E�  �        �� W�E� W        �E�  �        �E� W        P�a� �a�e� Q        ]�d� r        ��� R���� �        ��� q        ��� r  ����� R        ��ǩ � ǩש P        ���� ����� Rǩש R        ��ǩ J�        ��Ʃ SƩǩ � � <"�        ��ũ s        ��ǩ 	��        ��Ʃ s�Ʃǩ � � <"#�        ��ǩ Q        ���� s	����© R©ũ s	��        �� ��� Q        �� � � <"��� � r "�        �� � � <"#         �� ��� Q        �� � � <"��� � r "�        �� � � <"#        p�x� Qx��� uT��� uT߫� Q�l� uT���� uT�� Q�� uTC�X� QX�o� uTq�u� Qu�v� uT{��� uT        U��� ���l� ����o� ��q��� ��        U�x� w߫� r�� rC�T� rq�u� r        �+� u        �߫ S��� S�C� Sv�{� S���� S        5�<� P        #�+� u        #�1� P        :�T� S        D�T� 1�        D�P� R        D�K� r        ���� v����� V        u�߫ S��� S�C� Sv�{� S���� S        ��߫ uT        u��� W��ά Rά� W�*� R*�C� Wv�z� Rz�{� W���� W        ���  ��C�  �v�{�  �����  �        ��ά Rά� W�*� R*�C� Wv�z� Rz�{� W���� W        ��ˬ Pˬά r� �*� P*�A� uTv�z� Pz�{� uT���� uT        ���  ��C�  �����  �        ��ˬ Pˬά r� �*� P*�A� uT���� uT        �C�  �����  �        �A� uT���� uT        ���� uT��߫ uT        ���� P��ͫ P        ī߫ uT        īͫ P        ī߫ ��           ѫث P        ���� 1�        ֫߫ S        �� uLu��� v��&� V���� V�� uLu�C�o� uLu�q�v� uLu�{��� uLu�        �l� S���� S�� SC�o� Sq�v� S{��� S        �l� W���� W        �� R�� uP�� R�� uPC�X� RX�o� uPq�u� Ru�v� uP{��� uP        ��  �C�o�  �q�v�  �{���  �        �� R�� uPC�X� RX�o� uPq�u� Ru�v� uP{��� uP        ��� WC�m� Wq�v� W{��� W        ���  �C�o�  �{���  �        ��� WC�m� W{��� W        C�o�  �{���  �        C�m� W{��� W        �&� W*�l� W���� W        �� P*�=� P        2�l� W        2�=� P        2�l� �           A�H� P        �� 1�        F�l� S        P�l� 1�        P�\� R        P�W� r        ɪ� u        ɪ� u        ɪ� S        �� P        ٪� u        ٪� u        ٪� P        ��� R��� S        ��� 1�        ��� R        ���� r        ���� R        ���� 0�        ���� r        ��ŭ 1���� 1�        ��ŭ S�� S��� S        ��ŭ s��� s���� s�        ���� s        ح� 1�� � 1�        ح� V� � V        ح� v�� � v�        حܭ v        ��Ȫ u`�Ȫɪ t\�l��� u`����� t\�        ���� P        {��� 1�        {��� P        {��� p        K�Q� PQ�Z� p Z�_� �o        k�q� Pq�z� p z�� �o        ���� S���� �        ��Ѯ VѮҮ P        ��Ʈ R        ���� r        �� S�� ��0� S0�2� �        �� V�� P�1� V1�2� �         �� S�� �        �1� V1�2� P        �&� R        �!� r        M�n� Sn�p� �p��� S���� �        M�o� Vo�p� Pp��� V���� �         Q�n� Sn�p� �        p��� V���� P        z��� R        z��� r        ��� 0��*� 1�e��� 0�հ.� 0�2�\� 0�p��� 0�        ԯ*� We��� Wհ"� W)�.� W        ̯*� We��� Wհ.� W2�\� Wp��� W        ԯ� Se��� Sհ"� S)�.� S        e���  �հ"�  �)�.�  �        e��� Sհ"� S)�.� S        x��� P���� s� ���� uHհ� P�"� uH)�-� P-�.� uH        ~���  �հ"�  �        ~��� P���� s� ���� uHհ� P�"� uH        հ"�  �        հ"� uH        �*� V        ��� u���� t ���� t���� t���� t��� t�� t�� t        �*� S        ��� P�R�        �*� W        �*� 1�        �&� R        �!� r        H�\� 1�p�y� 1�        H�\� Vp�y� V        H�\� v�p�y� v�        H�L� v        ���� w        *�d� u`�d�e� t\���԰ u`�԰հ t\�        J�R� P        ��հ 1�        ��ǰ P        ��° p        ��� � �� R��� R        ��� ���� �        ı� � � <"#��� r r <"#        /��� 0����� 1�ղ� 0�E��� 0���̳ 0��� 0�        D��� Wղ� WE��� W���� W        <��� Wղ� WE��� W��̳ W��� W        D�U� Sղ� SE��� S���� S        ղ�  �E���  �����  �        ղ� SE��� S���� S        ��� P�� � s�  �� uHE�Z� PZ��� uH���� P���� uH        ��  �E���  �        ��� P�� � s�  �� uHE�Z� PZ��� uH        E���  �        E��� uH        U��� V        c�i� ui�l� t l�m� tm�n� tn�o� to�s� ts�t� tt�v� t        c��� S        n�r� P�R�        X��� W        ���� 1�        ���� R        ���� r        ��̳ 1��� 1�        ��̳ V�� V        ��̳ v��� v�        ���� v        �� � w        ��Բ u`�Բղ t\��D� u`�D�E� t\�        ��² P        +�E� 1�        +�7� P        +�2� p        0�9� �9�=� P        u�մ 0�մ� 1�*�c� 0���� 0��� 0�0�n� 0�        ��� V*�c� V��� V�� V        ��� V*�c� V��n� V        ���� W*�c� W��� W�� W        *�c�  ����  ���  �        *�c� W��� W�� W        8�M� PM�P� w� P�c� uH���� P��� uH�� P�� uH        >�c�  ����  �        >�M� PM�P� w� P�c� uH���� P��� uH        ���  �        ��� uH        ��� uD        ��˴ Q        ��� V        ��� S        ߴ� 1�        ߴ� R        ߴ� r        �� 1�0�9� 1�        �� S0�2� S4�9� S        �� s�0�2� s�4�9� s�        �� s        L�Z� Q`�d� Q        L�Z� q�`�d� q�        L�P� q        �)� u`�)�*� t\�c��� u`����� t\�        �� P        {��� 1�        {��� P        {��� p        p�y� �y�}� P        ���� 0���� 1�Q��� 0�ŷ� 0�"�L� 0�`��� 0�        ��� WQ��� Wŷ� W�� W        ��� WQ��� Wŷ� W"�L� W`�z� W        ��Ѷ SQ��� Sŷ� S�� S        Q���  �ŷ�  ���  �        Q��� Sŷ� S�� S        h�}� P}��� s� ���� u@ŷڷ Pڷ� u@�� P�� u@        n���  �ŷ�  �        n�}� P}��� s� ���� u@ŷڷ Pڷ� u@        ŷ�  �        ŷ� u@        Ѷ� V        ߶� uH        ߶� S        �� P�R�        Զ� W        �� 1�        �� R        �� r        8�L� 1�`�i� 1�        8�L� V`�i� V        8�L� v�`�i� v�        8�<� v        |��� w        �P� u`�P�Q� t\���ķ u`�ķŷ t\�        6�>� P        ��ŷ 1�        ���� P        ���� p        ۸,� 0�,�F� 1���ù 0���N� 0�R�|� 0���κ 0�        �F� W��ù W��B� WI�N� W        �F� W��ù W��N� WR�|� W���� W        �� S���� S��B� SI�N� S        ��ù  ���B�  �I�N�  �        ���� S��B� SI�N� S        ���� P���� s� ��ù u@��
� P
�B� u@I�M� PM�N� u@        ��ù  ���B�  �        ���� P���� s� ��ù u@��
� P
�B� u@        ��B�  �        ��B� u@        �F� V        �F� uH        �F� S        �� P�R�        �F� W        6�F� 1�        6�B� R        6�=� r        h�|� 1����� 1�        h�|� V���� V        h�|� v����� v�        h�l� v        ���� w        F��� u`����� t\�ù�� u`����� t\�        f�n� P        ۹�� 1�        ۹� P        ۹� p        �V� 0�V�p� 1���� 0��n� 0�r��� 0���� 0�        �p� W��� W�b� Wi�n� W        �p� W��� W�n� Wr��� W��ʼ W        �+� S��ܻ S�b� Si�n� S        ���  ��b�  �i�n�  �        ��ܻ S�b� Si�n� S        ��ͻ Pͻл s� л� u@�*� P*�b� u@i�m� Pm�n� u@        ���  ��b�  �        ��ͻ Pͻл s� л� u@�*� P*�b� u@        �b�  �        �b� u@        +�p� V        9�p� uH        9�p� S        D�H� P�R�        .�p� W        `�p� 1�        `�l� R        `�g� r        ���� 1����� 1�        ���� V���� V        ���� v����� v�        ���� v        ̼м w        p��� u`����� t\��� u`��� t\�        ���� P        ��� 1�        ��� P        ��� p        ?��� 0����� 1��#� 0�U��� 0���ܾ 0��.� 0�        T��� W�#� WU��� W���� W        L��� W�#� WU��� W��ܾ W�
� W        T�e� S�� SU��� S���� S        �#�  �U���  �����  �        �� SU��� S���� S        ��� P�� s� �#� uHU�j� Pj��� uH���� P���� uH        ��#�  �U���  �        ��� P�� s� �#� uHU�j� Pj��� uH        U���  �        U��� uH        e��� V        s�y� u        s��� S        ���� P�R�        h��� W        ���� 1�        ���� R        ���� r        Ⱦܾ 1���� 1�        Ⱦܾ V��� V        Ⱦܾ v���� v�        Ⱦ̾ v        �� w        ��� u`��� t\�#�T� u`�T�U� t\�        нؽ P        ;�U� 1�        ;�G� P        ;�B� p        _��� 0���ʿ 1��C� 0�u��� 0����� 0��N� 0�        t�ʿ W�C� Wu��� W���� W        l�ʿ W�C� Wu��� W���� W�*� W        t��� S�<� Su��� S���� S        �C�  �u���  �����  �        �<� Su��� S���� S        �-� P-�0� s� 0�C� uHu��� P���� uH���� P���� uH        �C�  �u���  �        �-� P-�0� s� 0�C� uHu��� P���� uH        u���  �        u��� uH        ��ʿ V        ���� u���� t ���� t���� t���� t���� t���� t���� t        ��ʿ S        ���� P�R�        ��ʿ W        ��ʿ 1�        ��ƿ R        ���� r        ���� 1��� 1�        ���� V�� V        ���� v��� v�        ���� v        ,�0� w        ʿ� u`��� t\�C�t� u`�t�u� t\�        �� P        [�u� 1�        [�g� P        [�b� p        `�q� � q�u� pd�        d�q� � q�u� pd�        ���� S���� �         ���� P        �� P        �� S        �� P        0�;� �         v��� R        R��� S���� �         �� � v p "1� ��	 �p "1�         �7� � C�i� �          �;� �C�i� �        0�3� R3�7� �         0�B� P        C�Z� RZ�i� �         ���� �        ���� 0�        ���� V���� ����� V���� �        ���� 3�        ����
 ���������        ���� S���� P���� S���� �         )�@�
 v v <"�T�h� v p "����� v p "�        2�R� ST��� S        6��� :�        6�R� ST��� S        T��� :�        T��� S        ���� S���� �         �m� �m��� u���� t ��� u�:� WP�v� u���� u���� t���� u��� W�)� u7�_� W_�s� �s��� W���� u���� W���� W��� W        )�P� 0�P�d� Rd�g� r 4!�g�t� R���� R��� 0�        G�I� PI�:� uL��� uL        G�:� 	����� 	��        Y�b� Sb�:� uT��_� uT_�b� Sb�h� v v <"#xh�� uT        m��� P���� P���� P        D�_� ��Y  _�b� P	�� P�� w���� P���� w���� p����� P��� q�	� P_�s� ��Y          _�b� P        _�s� uT        ���� R��� S�7� S���� S        ��� ��Y  �7� ��Y  ���� ��Y          ���� R���� S        ���� W        ���� W        ���� t         ��� W�#� W#�7� uT���� uT        ��� S�7� S���� S        �� W�#� W#�7� uT���� uT        	�� P�� w        �7� uT���� W        ��� �TZ  7�_� �TZ  s��� �TZ  ���� �TZ          ��� Q�� uT7�K� QK�_� uTs��� uT���� uT        ��� 	��7�_� 	��s��� 	������ 	��        O�T� P���� P        ��� 1�        7�T� uT���� S���� uT        �� uTs��� uT        �	� P        s��� uT        ���� W���� W���� uT���� uT        ���� 1�        ���� uT���� W        $�:� 1���� 1�        $�:� S��� S        $�:� s���� s�        $�(� s        ���� 1����� 1�        ���� V���� V        ���� v����� v�        ���� v        d�g� 4�        d�g� �Z          q�t� R        q��� W        q�u� w        d�R� 0�]��� 0���C� 0�C�^� 2�f�� 0�        n��� S��R� uH]��� uH��f� uHf�z� Sz��� uH        n�R� 	��]��� 	����� 	��        |�� P��� W��R� uP]��� uP��f� uPf�i� Wi�o� uu<"#xo�� uP        ���� P�R� P]��� P���� PC�F� P        ���� uO�#� uOw��� 1�        d�R� �`  ]��� �`  ��� �`          ���� P        f�z� uP        ��#� V        ��#� �I`          ���� V        ���� S        
�#� uP        �#� S        ��#� uP        ���� uP�C� uP���� uP        ���� 	���C� 	������ 	��        .�6� P���� P        ���� 1�        �C� uP���� W        ���� uP        ���� S        ���� uP        	�� uPz�}� W}��� uP        �� 1�        z��� uP        Q�^� 2�        Q�]� R        Q�X� r        ���� 1���� 1�        ���� W��� W        ���� w���� w�        ���� w        ���� 1��� 1�        ���� W�� W        ���� w��� w�        ���� w         ��� ����� u���� u�J� S,�9� uD�|� S|��� ����� S���� ���� �         ��� 0����� uP���� uP���� uP��� uPY�e� uP�J� uPD�|� uP|��� 0����� uP���� 0����� uP��� 0��� uP         ��� 0����� 2���� 0�;�e� 0�g�� 0�        l�p� Rp�� u�;�� u�        |��� P���� uD;��� uD���� uD        ���� 	��;��� 	������ 	��        ���� P���� V���� uL;�|� uL|�� V��� uu<"#x���� uL���� uL        ���� P���� PJ�U� P        ���� P        |��� uL        v��� V,�3� V        -�t� Vg�� V��B� V��,� V        -�t� St�v� Vg�{� S{��� u@#���B� u@#���,� u@#�        -���  �g��  ���B�  ���D�  �        -��� uDg�� uD��B� uD��D� uD        g��� S��B� S��,� S        {��� s ���� W���� W�B� W��,� W        {���  ���B�  ���,�  �        {��� uD��B� uD��,� uD        {��� 0����� uT�B� uT��,� uT        {��� 0����� Q���� u����� Q���� q����� Q��1� Q1�B� u����� Q���� u����� Q���� u���� Q�,� u�        {��� 1����� P�1� P���� P���� P��� P�� 1q �$��� P        ���� P=�B� P���� P���� P'�,� P        v��� W        v�{� u~��� t         ���� W,�D� W        ���� V,�3� V        ���� P���� w        ,�D� uL        �J� uLD�G� VG�|� uL���� uL        �J� 	��D�|� 	������ 	��        S�`� P���� P        1�7� 1�        D�e� uL���� V���� uL        7�J� uLe�|� uL        ?�B� P        e�|� uL        ���� P��'� V�!� V!�&� P&�7� w J�U� PU��� VB��� VD�M� w         ����  �g�|�  �����  �����  �        ���� W���� uDg�J� uDJ�U� WU�|� uD���� uD���� uD        U��� SB��� S        c��� Q���� u@���� Q���� u@B�k� Qk�~� u@~��� Q���� u@���� Q���� u@        s��� P����
 1u@��$����� P����
 1u@��$�B�R� PR�Y� 1q �$�Y�k� Pk�~�
 1u@��$�~��� P����
 1u@��$����� P����
 1u@��$�        ���� P���� PR�Y� Pw�~� P���� P���� P        ���� ��e  g�|� ��e  ���� ��e  ���� ��e          ���� v pt"����� v r "�N�Y� w pt"�Y�\� w r "�        ���� 0�N�g� 0�        ���� v pt"#N�Y� w pt"#        ��� 1��� 1�        ��� V�� V        ��� v��� v�        ���� v        ���� 1�        ���� V        ���� v�        ���� v         �0� V         �'� v        #�@� 0�{��� 0��
� uT#�
�&� uTL�q� uT���� 0����� uT��� 0�        #�J� 0�{��� 0����� 2���J� 0�J�n� 2�n�x� 0�        ���� Q���� uL��� uL        ���� P���� uD        ���� 	��        ���� P���� V���� uH���� V���� uu<"#x���� uH        ��� P���� P5�J� Pn�u� P`�q� 	������ P        {��� u���� u��� u        ���� P        ���� uH        ���� v w ����� V        �&� uHL�O� VO�q� uH���� uH        �&� 	��L�q� 	������ 	��        [�q� P���� P        �� 1�        L�q� uH���� V        �&� uH        ���� P        &�J� uH        W��� V��� V�b� V��L� V        W��� S���� V�+� S+��� u@#��b� u@#���L� u@#�        W���  ����  ��b�  ���L�  �        W��� uD��� uD�b� uD��L� uD        ��� S�b� S��L� S        +�:� s :��� W�� W#�b� W��L� W        +���  ��b�  ���L�  �        +��� uD�b� uD��L� uD        +�:� 0�:��� uP#�b� uP��L� uP        +�:� 0�=�{� Q{��� u����� Q���� q����� Q�Q� QQ�b� u����� Q���� u���� Q�� u��;� Q;�L� u�        +�:� 1�I�{� P#�Q� P���� P��� P�"� P"�'� 1q �$�'�;� P        ���� P]�b� P���� P�� PG�L� P        ���� W        ���� V        ���� W        ��� V�� QL�W� Qq��� Q        ���� u        ��&� SL��� S���� S        ��� �tq  q��� �tq          ���� p r "�        ��� uL�U� uq��� u        ��&� SL��� S���� S        ��� pt�q��� pt�        q��� S        q��� pt�        ���� p s "�        �� P�Q� V��� V�� Qn�u� Pu�� Vb��� VL�W� Qq��� Q        �J�  �n���  �����  �        �� W�J� uDn�u� Wu��� uD���� uD        u�� Sb��� S        ���� Q���� u@���� Q��� u@b��� Q���� u@���� Q���� u@���� Q���� u@        ���� P����
 1u@��$����� P���
 1u@��$�b�r� Pr�y� 1q �$�y��� P����
 1u@��$����� P����
 1u@��$����� P����
 1u@��$�        ���� P	�� Pr�y� P���� P���� P���� P        ��J� �m  n��� �m  ���� �m          ���� w pt"����� w r "���� w pt"��� w r "�V�a� w pt"�a�c� w r "�        ���� 0���� 0�V�n� 0�        ���� w pt"#��� w pt"#V�a� w pt"#        ���� 1��-� 1�        ���� V�-� V        ���� v��-� v�        ���� v        D�R� Qc�g� Q        D�R� q�c�g� q�        D�H� q        V�f� W        V�]� w        ���� 0���� 0��#� w�#�5� Ws��� W���� w����� W���� 0����� W��� 0�n�y� Wy�{� 0�        ���� 0����� 0����� 0���n� 0�s��� 0�        ���� uH���� uH,�.� uHn�{� uH        ���� 	������ 	��,�.� 	��n�{� 	��        ���� S���� S,�.� Sn�{� S        �� P���� p ���I�X� P���� 	��        #�5� Ss��� Sn�y� S        #�5� 	��s��� 	��n�y� 	��        -�5� S        ���� P        5�X� S        ���� Pn�q� P        '�-� 1�        s��� Sn�y� S        E��� ��u          E�V� QV��� uT        E�V� RV��� uP        w��� S        ���� S        ��5� �v  s��� �v  n�y� �v          ���� 	��        ���� u        ���� Q��5� uTs��� uTn�y� uT        �� ��x  ���� ��x          �� p r "�        
�-� us��� u���� u        �5� uTs��� uTn�y� uT        �� pt����� pt�        ���� uT        ���� pt�        ���� p uT"�        ��� u���� u��� uy�{� u        ��
� ��u  
�� P���� P'�*� P*�-� s���� P���� s���� ��u  y�{� ��u          
�� P        ���� Sy�{� S        ���� S���� S        ���� 1�        ���� S        �,� 1�.�C� 1�        �,� W.�C� W        �,� w�.�C� w�        �!� w        Z�n� 1�{��� 1�        Z�n� S{��� S        Z�n� s�{��� s�        Z�^� s        ���� W        ���� w         �� ��� R�� r��!� R         �� �� � S �!� �         �� 0��� P�� P        X�l� Sl�p� �         ���� S���� �         ���� S���� �         ���� S�� � �         8�L� SL�P� �         h�|� S|��� �         ���� S���� �         ���� S�� � �         �,� S,�0� �         H�\� S\�`� �         x��� S���� �         H�\� S\�`� �         X�l� Sl�p� �         ���� P���� �P�        ���� R���� �R�        ���� p����� �P#�        ���� Q���� s�        ���� P���� S��o� uL�o�p� tH�p��� uL����� tH����� uL����� S����� uL�        �� P��o� uH�o�p� tD�p��� uH����� tD����� uH�        �G� Sp��� S���� S        �� Q�o� uPo�p� tLp��� uP���� tL���� uP        �� P�m� Vp��� V���� V        �� R�o� uTo�p� tPp��� uT���� tP���� uT        ���� ug����� P���� ug����� P��o� ug�o�p� tc�p��� ug����� tc����� ug�        ��� u���� u        ��� u���� u        ���� ug����� P��o� ug�o�p� tc�p��� ug����� tc����� ug�        ��� u���� u        ��� u���� u        �*� P|��� P���� S        "�0� S        0�:� V        L�p� �{)  ���� �{)          R�Y� ug����� ug�        R�\� P���� P        Y�p� �k)  ���� �k)          _�f� ug����� ug�        _�k� P���� P        ���� ug����� R���� ug�        ���� P���� uL<�        ���� P��� V�� �P��/� V/�0� �P�        ���� R��0� �R�        8�T� ST�V� uV�Z� t[�n� S        x��� S���� u���� t���� S        ���� S���� u���� t��� S        5�B� P�B�B� uH�B�E� �@�E�V� uH�V�Y� tD�]�y� uH����� uH�        5�B� PB�X� uHX�@� VE�T� V]�_� V���� V���� uH���� V���� V        E�O� RO�B� uLB�E� �DE�V� uLV�Y� tH]�y� uL���� uL        H�O� PO�� uT��B� uTB�E� �LE�V� uTV�Y� tP]�_� uT���� uT���� uT        X��� W���� 0����� P��A� WE�U� W]�_� W���� W���� 0����� 0�        +�4� P4�B� ug�B�E� �_�E�V� ug�V�Y� tc�Y��� ug�        +�:� V:�X� uY�[� V[�]� u���� u        +�U� WU�X� uY�]� W���� W        �X� uY�]� u���� u        +�.� s         m�{� P{��� p����� uT1����� P���� uT1����� uT1�        ���� V        ��� 0�        ���� Q��� uP        ��� �	1          ���� p r "�        ��� uP        ��� pt�        ��� uP        ��� pt�        �� p uP"�        )�Y� �\/          2�B� ug�B�E� �_�E�V� ug�V�Y� tc�        2�>� P>�B� uH<�B�E� �@<�E�L� PL�V� uH<�V�Y� tD<�        d�y� �\/          j�t� ug�t�x� Rx�y� ug�        j�x� Px�y� uH<�        ~��� ug����� R���� ug�        ~��� P        ��S� �S�c� p c��� �        ���� P        ��9� 0�9�@� P@��� W         �� P�� ��S�c� Pc��� ��        �� Pk�o� Po�~� S~��� P        ,�f� V        `��� U���� P��H� U        `��� W��H� W        i��� R���� 1w �$����� R��� 1w �$��*� R*�:� 1w �$�:�\� R\�l� 1w �$�l�x� Rx��� 1w �$����� R���� 1w �$����� R���� 1w �$����� R��� 1w �$��� R�(� 1w �$�(�8� R8�H� 1w �$�        ���� P�� P3�:� Pe�l� P���� P���� P���� P���� P���� P�� P!�(� PA�H� P        ]�~� R~��� u���� t���� u        ]��� S���� u���� t���� S        ���� R���� u���� t���� u        ���� S���� u���� t���� S        �� � R �*� u*�+� t+�>� u        ��(� S(�*� u*�+� t+�>� S        @�Y� � Y�a� Pa�b� �         Q�Y� �         p��� � ���� P���� �         ���� �         ���� P���� �        �$� P$�9� �        y��� P���� �        ���� P���� �         �8� � 8�A� PA�B� �         1�8� �         h�k� Rk�v� �        ���� R���� �        ��� R�(� u(�)� t)�<� u        ��&� S&�(� u(�)� t)�<� S        M�m� Rm�w� uw�x� tx��� u        M�u� Su�w� uw�x� tx��� S        ���� R���� u���� t���� u        ���� S���� u���� t���� S        ���� � ��� P�� �         ���� �         �)� � )�1� P1�2� �         !�)� �         Y�d� Pd�y� �        ���� P���� �        �$� P$�9� �        y��� P���� �        ���� � ���� P���� �         ���� �         �� R�� �        X�[� R[�f� �        ���� �V�Z� �k�|� �        ���� R��� u�� t�Q� uQ�R� tR�|� u        ��� S�� u�� t�N� SN�Q� uQ�R� tR�|� S        ���� �&�*� �;�L� �        ���� R���� u���� t��!� u!�"� t"�L� u        ���� S���� u���� t��� S�!� u!�"� t"�L� S        ���� R���� u���� t���� u        ���� S���� u���� t���� S        ��� R�� u�� t�)� u        ��� S�� u�� t�)� S        =�]� R]�g� ug�h� th�{� u        =�e� Se�g� ug�h� th�{� S        ���� � ���� P���� �         ���� �         ���� � ���� P���� �         ���� �         ��� P�� �        Y�d� Pd�y� �        ���� P���� �        `��� ��� ��)� �        q��� Q���� u���� t���� u���� t��)� u        q��� S���� u���� t���� S���� u���� t��)� S        ���� R���� u���� t��� u        ���� S���� u���� t��� S        �5� R5�M� uM�N� tN�a� u        �K� SK�M� uM�N� tN�a� S        ���� R���� u���� t��J� u        ���� S��J� S        ���� P���� ud�� ud        ���� P��� ud        ���� ����� � ##(        o� R�� �        o� S�� � �� S        �� R�� �        �� S�� � �� S        Z] �         `� �        � �        �� R�� �        �� S�� � �� S        �� ��� p �� �        �� R�� �        �� S�� �         @| ��� ��� �        Qc Rc� u�� t�� u�� t�� u        Q� S�� u�� t�� S�� u�� t�� S        �	 P        	&	 Q2	6	 Q        @	�	 �[
`
 �        @	n	 �n	�	 U�		
 W	
m
 U�
�
 W�
 U\ W\z Uz� W�� U        n	�	 V        e	h	 Ph	� �        �	�	 0��	
 S�
�
 S\ 0�z� 0��� S        �	
 S�
�
 SKW SW\ R�� S        �	`
 0��
�
 0�\ 0�z� 0�        �	�	 R- Rz� R�� �P        �	`
 V�
�
 V\ Vz� V        -K P        �	
 0��
�
 0��� 0�        �	
 U�
�
 U�� U        �	
 V�
�
 V�� V        �
�
 P        �	m
 0��
� 0�        �	�	 S�
 S\z S�� S        �	m
 V�
� V         P        �
�
 P�� P        �
�
 �d  �� �d          �
�
 P�� P        �
�
 �H�� W        �
�
 1�        �� P        5I PI �P        `� S�8 SAU RU� S� R S        `_ �Ld �L        `� U� U        Ad �g  � �g          CZ V� V        OU 1�        � V        `q 	��q W�� 	���� W<I 	��IU PUm 	���� W
 P        �� V<U V
 V        �� WIU P
 P        �� P        <U V
 V        IU P
 P        � �$g �� �g �� �Fk  d� �$g �� �Xj  �� �g �� �Fk  |� �$g �� �Xj  �� �g �� �Fk          q �"i  � �Nj  �� �$j  �� �$j  �� �<k  d� �Nj  �� �<k  Um �"i  |� �Nj  �� �<k  �
 �$j          q� �$g  �< �$g  U
 �$g          q� 	���< 	��U
 	��        q� 	���� �Td� 	���� �TUm 	��|� 	���� P�� �T        d� �X|� Q�� �X        �� �T�� P�� �T        �� P�� �X#        �� �X        �� P�� �T        5 R        �� �g  �� �g  �� �g  �
 �g          �� 	���� 	���� 	���
 	��        �� 	���� W�� 	���� W�� 	���� P�� W�
 	��        �� V�� V        �� W�� W�� P�� W        �� P        �� V        �� P�� W        �d *��< *�        � P�� P2 P        �d �P�< �P        �� P        $ P$8 u s �        m| 4�        m| �,        mw �,         / �/3 V���3� V�W��� V�W��B V�W�Ts V�W�         � ��1 �        7� U�� ��� U�x �        �� ��l  �x ��l          �� �l  �x �l          �� 	���x 	��        �� 	���� W�� 	���� W1i 	��ix P        �� VTx V        �� Wix P        �� P        �� ��l � ��l  �o   ��l 1 �o          �� ��m  �� �
o  �� ��n  �1 �
o  1T ��m          �� ��l  �T ��l          �� 	���T 	��        �� 	��� 	�� 	��/ P1T 	��        �1 �        / P        1 �        �� 2�        �� �        �� �        �� 4�        �� �        �� �        �� P        �� Q�� Q        �� P        � Q Q        -A P        <V Qbf Q        �� P�� V'� V�� V)E VIS VU] Vkr V�� V        �� 0��� u@�� t��& u@&' t�'� u@�� 0��v u@v� 0��� u@�� 0��� u@)E u@I] u@k� u@        �� 0��� u��� t��& u�&' t�'� u��� 0��� u�� 0�- u�-@ 0�@M u�M� 0��� 0�)E 0�I] u�k� u�        �P 0�P� u��� t��& u�&' t�'B u�Be 0�e� u��  0� - u�-� 0��� 0�)E 0�IM 0�MQ u�QS 0�SU u�U] 0�kr 0�r� u��� 0�        �� uD�� t@�& uD&' t@        �� V        �� uP��� tL��& uP�&' tL�'� uP��� uP��� uP��E uP�I] uP�k� uP�        �� uP��� tL��& uP�&' tL�'� uP��� uP��� uP��E uP�I] uP�k� uP�        �� ud��� t`��& ud�&' t`�'� ud��� ud��� ud��E ud�I] ud�k� ud�        �� Q�� uDv� Q�� uD        v� ud��� P�� ud�        v� uD        v� 	��        v� uD#�        �� W        �� V'� V�v V�� V�� V)E VIS VU] Vkr V�� V        � V        #� uT��� tP��& uT�&' tP�'� uT��v uT�I] uT�k� uT�        &� ud��� t`��& ud�&' t`�'� ud��v ud�I] ud�k� ud�        &2 RMm R        Md ud�dm Pmv ud�        Mm R        Mv 	��        Mm r�        Sm Qmv w�        U� V'� V�M VIS VU] Vkr V�� V        e~ V        ~� uX��� tT��& uX�&' tT�'� uX��� uX�M uX�I] uX�k� uX�        �� uX��� tT��& uX�&' tT�'� uX��� uX�M uX�I] uX�k� uX�        �� ud��� t`��& ud�&' t`�'� ud��� ud�M ud�I] ud�k� ud�        �� P-7 P        �� V'� V�� V- V@M VIS VU] Vkr V�� V        �� VIK V        �� u\��� tX��& u\�&' tX�'� u\�- u\�@M u\�KQ u\�SY u\��� u\�        �� ud��� t`��& ud�&' t`�'� ud�- ud�@M ud�KQ ud�SY ud��� ud�        �� P@G P        �� V'� V- VKQ VUY V�� V        ' VWY V�� V        '� u`��� t\��& u`�&' t\�'B u`�e� u`�- u`�KQ u`�SU u`��� u`��� u`�        8� u`��� t\��& u`�&' t\�'B u`�e� u`�- u`�KQ u`�SU u`��� u`��� u`�        8� ud��� t`��& ud�&' t`�'B ud�e� ud�- ud�KQ ud�SU ud��� ud��� ud�        8> P P        S� V'B Ve� V - VMQ V�� V        c| V        �� ud��� t`��& ud�&' t`�e� ud� - ud�        �� u`��� t\��& u`�&' t\�e� u`� - u`�        �� P ' P        �� Ve� V        �� V        �� Ve~ V        �� V        �P WP� s&��� w\��� W�# s&�#% w\�        �V v$��� v$�        �V V�� V        �� uD�� t@�& uD&' t@        J W        J v$�        J V        J uD        V� W�% W        V� v��$ v�        V� V�$ V        V� uD�� t@�& uD&' t@        y� W        y� v�        y� V        y� uD�� t@        �� uT�        �� ud��� R�� ud�        �� P        �� ud�        �� u`�        �� P        �� ud��� R�� ud�        �� P        �� P        �� Q Q        1 P        ,F QRV Q        m� P        |� Q�� Q        �� P�  S�� S�� S7< SVZ S\^ S�� S�� S�� S�� S 7  S        j 0�jX u�XY t�Y� u��� t��� u��� 0�m u�m� 0��� u�3 u�7H u�V� u��� 0��� u��� 0��7  u�        - 0�-X u�XY t�Y� u��� t��r u�r� 0�  0� m u�m� 0��� u��� 0��� u�3 u�7< 0�<H u�VX u�X\ 0�\^ u�^� 0��+  u�+ -  0�- 2  u�2 7  0�        � 0��X u�XY t�Y� u��� t��2 u�2� 0�- 0�-M u�M` 0�`m u�m� 0��� u��� 0��� u�3 0�7< 0�<H u�V� 0��  u�   0� $  u�$ 7  0�        | 0�|X u�XY t�Y� u��� t��� u��� 0�@ 0�@M u�M� 0��� u�3 0�7H 0�V� 0��� u��� 0��� u��7  0�        �� S        �  S�� S� S�� S7< SVZ S\^ S�� S�� S�� S�� S 7  S        �� S          S�� S� S�� S7< SVZ S\^ S�� S�� S�� S�� S 7  S         S        X u�XY t�Y� u��� t�          S�� S� S�� S7< SVZ S\^ S�� S�� S�� S�� S 7  S        (A S        AX uH�XY tD�Y� uH��� tD��� uH� uH�3 uH�7H uH�V� uH��� uH��7  uH�        RX uH�XY tD�Y� uH��� tD��� uH� uH�3 uH�7H uH�V� uH��� uH��7  uH�        RX ud�XY t`�Y� ud��� t`��� ud� ud�3 ud�7H ud�V� ud��� ud��7  ud�        RX Pmw P        m  S�� Sm S�� S�� S7< SVZ S\^ S�� S�� S�� S�� S�� S�� S 7  S        }� S�� S�� S        �X uL�XY tH�Y� uL��� tH��� uL�m uL��� uL��� uL�3 uL�7H uL�VX uL�\^ uL��7  uL�        �X ud�XY t`�Y� ud��� t`��� ud�m ud��� ud��� ud�3 ud�7H ud�VX ud�\^ ud��7  ud�        �� P�� P        �  S�� Sm S�� S7< SVX S\^ S�� S�� S�� S�� S 7  S        � S�� S7< S        X uP�XY tL�Y� uP��� tL��r uP�m uP��� uP�3 uP�<H uP�VX uP�\^ uP��+  uP�- 2  uP�        X uP�XY tL�Y� uP��� tL��r uP�m uP��� uP�3 uP�<H uP�VX uP�\^ uP��+  uP�- 2  uP�        X ud�XY t`�Y� ud��� t`��r ud�m ud��� ud�3 ud�<H ud�VX ud�\^ ud��+  ud�- 2  ud�         P P        0  S�r S m S�� SVX S\^ S�� S�� S�� S�� S +  S- 2  S        @Y SVX S\^ S        mX uT�XY tP�Y� uT��� tP��R uT� m uT��� uT�<H uT��)  uT�        pX ud�XY t`�Y� ud��� t`��R ud� m ud��� ud�<H ud��)  ud�        p{ P ' P        �  S�R S-m S�� S�� S�� S�� S�� S )  S        �� S�� S�� S        �X uX�XY tT�Y� uX��� tT��2 uX�-m uX��� uX�<H uX��� uX��� uX��  uX� $  uX�        �X uX�XY tT�Y� uX��� tT��2 uX�-m uX��� uX�<H uX��� uX��� uX��  uX� $  uX�        �X ud�XY t`�Y� ud��� t`��2 ud�-m ud��� ud�<H ud��� ud��� ud��  ud� $  ud�        �� PMW P        �  S�2 S-M S`m S�� S�� S�� S�� S�� S   S $  S        �� S�� S   S        X u\�XY tX�Y� u\��� tX�� u\�-M u\�`m u\��� u\��� u\��� u\�   u\�        X ud�XY t`�Y� ud��� t`�� ud�-M ud�`m ud��� ud��� ud��� ud�   ud�        ! P`g P        '  S� S-M S�� S�� S�� S�� S   S        7S S�� S        SX u`�XY t\�Y� u`��� t\��� u`�-M u`��� u`�        dX u`�XY t\�Y� u`��� t\��� u`�-M u`��� u`�        dX ud�XY t`�Y� ud��� t`��� ud�-M ud��� ud�        dj P-7 P          S�� S@M S�� S        �� S        �X ud�XY t`�Y� ud��� t`��� ud�@M ud�        �X u`�XY t\�Y� u`��� t\��� u`�@M u`�        �� P@G P        �  S�� S        �� S        �  S�� S        �� S         W WY� W         U s�Y� s�         U SY� S         X u�XY t�Y� u��� t�        7W W        7U s�        7U S        7X u�XY t�        # uT�         ud�  R # ud�          P        ^� uL�        dn ud�nr Rr� ud�        dr P        �� ud�        �� u`�        �� P        �  u\�        �  ud� 	  R	   ud�        �	  P        M a  P        \ v  Q� �  Q        � �  P�  $ Ss$}& S&�& S'' S6':' S<'>' Sy'�' S�'�' S�'�' S�'�' S�'( S        � J! 0�J!8$ u�8$9$ t�9$r$ u�r$s$ t�s$�% u��%�% 0��%M& u�M&`& 0�`&�& u��&' u�'(' u�6'{' u�{'}' 0�}'�' u��'�' 0��'( u�        � " 0�"8$ u�8$9$ t�9$r$ u�r$s$ t�s$R% u�R%�% 0��% & 0� &M& u�M&v& 0�v&& u�&�& 0��&�& u��&' u�'' 0�'(' u�6'8' u�8'<' 0�<'>' u�>'�' 0��'( u�(( 0�(( u�(( 0�        � �" 0��"8$ u�8$9$ t�9$r$ u�r$s$ t�s$% u�%�% 0��%& 0�&-& u�-&@& 0�@&M& u�M&v& 0�v&{& u�{&�& 0��&�& u��&' 0�'' 0�'(' u�6'�' 0��'�' u��'�' 0��'( u�(( 0�        � \# 0�\#8$ u�8$9$ t�9$r$ u�r$s$ t�s$�$ u��$�% 0��% & 0� &-& u�-&�& 0��&�& u��&' 0�'(' 0�6'�' 0��'�' u��'�' 0��'�' u��'( 0�        � �  S        �  $ Ss$�% S�%}& S&�& S'' S6':' S<'>' Sy'�' S�'�' S�'�' S�'�' S�'( S        � �  S        �  $ Ss$�% S�%}& S&�& S'' S6':' S<'>' Sy'�' S�'�' S�'�' S�'�' S�'( S        � �  S        �#8$ u�8$9$ t�9$r$ u�r$s$ t�        �  $ Ss$�% S�%}& S&�& S'' S6':' S<'>' Sy'�' S�'�' S�'�' S�'�' S�'( S        !!! S        !!8$ uH�8$9$ tD�9$r$ uH�r$s$ tD�s$�% uH��%�& uH��&' uH�'(' uH�6'{' uH�}'�' uH��'( uH�        2!8$ uH�8$9$ tD�9$r$ uH�r$s$ tD�s$�% uH��%�& uH��&' uH�'(' uH�6'{' uH�}'�' uH��'( uH�        2!8$ ud�8$9$ t`�9$r$ ud�r$s$ t`�s$�% ud��%�& ud��&' ud�'(' ud�6'{' ud�}'�' ud��'( ud�        2!8! PM&W& P        M! $ Ss$�% S�%M& S`&}& S&�& S'' S6':' S<'>' Sy'{' S}'�' S�'�' S�'�' S�'�' S�'�' S�'( S        ]!v! Sy'{' S}'�' S        �!8$ uL�8$9$ tH�9$r$ uL�r$s$ tH�s$r% uL��%M& uL�`&m& uL�o&& uL��&' uL�'(' uL�6'8' uL�<'>' uL��'( uL�        �!8$ ud�8$9$ t`�9$r$ ud�r$s$ t`�s$r% ud��%M& ud�`&m& ud�o&& ud��&' ud�'(' ud�6'8' ud�<'>' ud��'( ud�        �!�! P`&g& P        �! $ Ss$r% S�%M& So&}& S'' S6'8' S<'>' S�'�' S�'�' S�'�' S�'�' S�'( S        �!�! So&t& S'' S        �!8$ uP�8$9$ tL�9$r$ uP�r$s$ tL�s$R% uP��%M& uP�t&& uP��&' uP�'(' uP�6'8' uP�<'>' uP��'( uP�(( uP�        �!8$ uP�8$9$ tL�9$r$ uP�r$s$ tL�s$R% uP��%M& uP�t&& uP��&' uP�'(' uP�6'8' uP�<'>' uP��'( uP�(( uP�        �!8$ ud�8$9$ t`�9$r$ ud�r$s$ t`�s$R% ud��%M& ud�t&& ud��&' ud�'(' ud�6'8' ud�<'>' ud��'( ud�(( ud�        �!�! P�%�% P        " $ Ss$R% S &M& Sv&}& S6'8' S<'>' S�'�' S�'�' S�'�' S�'�' S�'( S(( S         "9" S6'8' S<'>' S        M"8$ uT�8$9$ tP�9$r$ uT�r$s$ tP�s$2% uT� &M& uT�v&{& uT�'(' uT��'	( uT�        P"8$ ud�8$9$ t`�9$r$ ud�r$s$ t`�s$2% ud� &M& ud�v&{& ud�'(' ud��'	( ud�        P"[" P && P        a" $ Ss$2% S&M& Sv&{& S�'�' S�'�' S�'�' S�'�' S�'	( S        q"�" S�'�' S�'�' S        �"8$ uX�8$9$ tT�9$r$ uX�r$s$ tT�s$% uX�&M& uX�v&{& uX�'(' uX��'�' uX��'�' uX��'�' uX��'( uX�        �"8$ uX�8$9$ tT�9$r$ uX�r$s$ tT�s$% uX�&M& uX�v&{& uX�'(' uX��'�' uX��'�' uX��'�' uX��'( uX�        �"8$ ud�8$9$ t`�9$r$ ud�r$s$ t`�s$% ud�&M& ud�v&{& ud�'(' ud��'�' ud��'�' ud��'�' ud��'( ud�        �"�" P-&7& P        �" $ Ss$% S&-& S@&M& Sv&{& S�'�' S�'�' S�'�' S�'�' S�'�' S�'( S        �"�" S�'�' S�'�' S        �"8$ u\�8$9$ tX�9$r$ u\�r$s$ tX�s$�$ u\�&-& u\�@&M& u\�v&{& u\��'�' u\��'�' u\��'�' u\�        �"8$ ud�8$9$ t`�9$r$ ud�r$s$ t`�s$�$ ud�&-& ud�@&M& ud�v&{& ud��'�' ud��'�' ud��'�' ud�        �"# P@&G& P        # $ Ss$�$ S&-& Sv&{& S�'�' S�'�' S�'�' S�'�' S        #3# Sv&{& S        3#8$ u`�8$9$ t\�9$r$ u`�r$s$ t\�s$�$ u`�&-& u`��'�' u`�        D#8$ u`�8$9$ t\�9$r$ u`�r$s$ t\�s$�$ u`�&-& u`��'�' u`�        D#8$ ud�8$9$ t`�9$r$ ud�r$s$ t`�s$�$ ud�&-& ud��'�' ud�        D#J# P&& P        _# $ Ss$�$ S &-& S�'�' S        o#�# S        �#8$ ud�8$9$ t`�9$r$ ud�r$s$ t`�s$�$ ud� &-& ud�        �#8$ u`�8$9$ t\�9$r$ u`�r$s$ t\�s$�$ u`� &-& u`�        �#�# P &'& P        �# $ Ss$�$ S        �#�# S        �# $ Ss$�$ S        �#�# S         $7$ W9$q$ W         $5$ s�9$o$ s�         $5$ S9$o$ S         $8$ u�8$9$ t�9$r$ u�r$s$ t�        $7$ W        $5$ s�        $5$ S        $8$ u�8$9$ t�        �&' uT�        �&�& ud��& ' R '' ud�        �& ' P        >'y' uL�        D'N' ud�N'R' RR'y' ud�        D'R' P        �'�' ud�        �'�' u`�        �'�' P        �'�' u\�        �'�' ud��'�' R�'�' ud�        �'�' P        -(A( P        <(V( Qb(f( Q        }(�( P        �(�( Q�(�( Q        �(�( P        �(�( Q)) Q        )") �").) S�P��)�) S�R�        H)I) PI)�) V9*�* V        ])g) PY*n* Pn*�* u�~        )�) u9*�* u        ])�) V9*�* V        �)5* W5*6* u�~�6*9* t�~�        �)4* V        �)6* u�~�6*9* t�~�        �)* S�R��**
 S�u�~��*3*
 S�u�~��3*6* p �u�~��6*9* p �t�~��        �)9* �S�          �)* V        �)* u�~�        �)* S        �*�* P        �*�* Q�*�* Q        +!+ P        +6+ QB+F+ Q        ]+q+ P        l+�+ Q�+�+ Q        �+�+ P�+�+ Q        �+�+ S         ,, P,+, Q        ,8, S        P,T, PT,{, Q        a,�, S        �,�, P�,�, Q        �,�, S        �,�, P�,- Q        -(- S        @-D- PD-k- Q        Q-x- S        �-�- P�-�- Q        �-�- S        �-�- P�-. Q        �-. S        0.4. P4.[. Q        A.h. S        �.�. P�.�. Q        �.�. S        �.�. P�.�. Q        �./ S         /$/ P$/K/ Q        1/X/ S        p/t/ Pt/�/ Q        �/�/ S        �/=0 � =0E0 PE0o0 Wu0�0 P�0�0 U�0�0 p v "#��0�0 p v "#��0�0 P�01 W11 p s "#�1&1 p s "#�&161 P61H1 � H1L1 WL1S1 U        �/E0 �E0S0 VS0Z0 v�Z0c0 Vu0�0 R�0�0 r v "#��0�0 r v "��01 R11 r s "#�1#1 r s "�#161 R61H1 �H1S1 R        �/�/ ��/u0 R61H1 R        �/�/ 0��/u0 Qu0�0 �h�01 Q1#1 U#1L1 QL1S1 �h        �/�/ 0��/�0 S�0�0 s��0�0 S61H1 SL1S1 S        �0�0 W�0�0 Q�0�0 �dL1S1 Q        �0�0 S�01 �q "H1L1 S        �1�1 W�1�1 ����1�1 v         �1�1 P�1�1 P        �1�1 Q�1�1 P�1�1 P        �1�1 r w ��1�1 R        �1�1 S�1�1 �        �1�1 P        +2-2 P        @2L2 �O2R2 P�u�        ~2�2 P�23 u@�56 u@�8�9 u@�9�9 u@*:^: u@        �23 W�5�5 W�5�5 w��56 W66 R6�6 u��7�8 u�        �2�2 V�2�2 uT#�5�5 q$�5 6 uT#$        �5�5 q(�5 6 uT#(        3T4 Vh4�4 V5:5 RA5�5 u@O7�7 V�8�8 R�9�9 R�9�9 u@�9�9 S�9�9 V�9�9 V        e203 u�5�6 u�7�8 u�8�9 u�9�9 u*:Y: uY:^: uDl�        ~2�2 uD�5�5 uD�8�9 uD�9�9 uD*:^: uD        �2�2 P�2�2 W�8�9 W�9�9 W*:^: W        �2�2 u#l#�8�8 u#l#        �8j9 0�j9�9 S�9�9 0��9�9 S*:3: 0�;:N: S        �8�9 0��9�9 0�;:N: 0�        �8�9 S�9�9 S;:N: S        �203 u �5�6 u �7�8 u         �23 S�5�5 S�56 S6�6 W�7$8 W.8�8 W        �2�2 W�23 P�5�5 P�56 W66 R6�6 u��7�8 u�        �2�5 8��5�5 8��5�8 8��9�9 8��9*: 8�        �23 u@�5�5 u@�56 u@         66 W66 R6�6 S�7)8 S.8�8 S        606 s 06�6 uT�6�6 u@�#0��7'8 uT'8.8 u@�#0�.8�8 uT        6�6 8��7�8 8�        606 0�06�6 V�6�6 P�6�6 V�78 V88 P8!8 V.8�8 V        606 0�36�6 Q�6�6 u��6�6 Q�7�7 Q�78 u�8=8 Q=8P8 u�P8]8 Q]8p8 u�p8}8 Q}8�8 u��8�8 Q�8�8 u��8�8 Q�8�8 u�        606 1�?6�6 P�7�7 P�7�7 1q �$��7�7 P�7�7 1q �$��7�7 P.8=8 PP8]8 Pp8}8 P�8�8 P�8�8 P        �6�6 P�7�7 P�7�7 P�78 PI8P8 Pi8p8 P�8�8 P�8�8 P�8�8 P        G3X3 RX3�3 S�3�4 u@O7[7 u@[7~7 S~7�7 u@�9�9 u@        �4�4 P�4�4 Q�4A5 u@�6O7 u@�8�8 u@�9�9 u@        �4�4 R�4�5 u��6O7 u��8�8 u��9�9 u�        3/3 u\�/343 P43s3 u\�s3z3 Pz3�3 u\��3�3 P�3�5 u\��6�7 u\��8�8 u\��9�9 u\��9*: u\�        +3/3 u\/303 p �4�4 w         3/3 u\�/343 P43s3 u\�s3z3 Pz3�3 u\��3�3 P�3r4 u\�r4u4 u`�u4�5 W�6O7 WO7�7 u\��8�8 W�9�9 W�9�9 u\��9�9 u\��9: W        �3�3 S        `34 0��9�9 0�        `3g3 s 1$�g3m3 Pm3p3 t p3u3 tu3v3 tv3z3 tz3�3 s 1$��34 u@1$��9�9 u@1$�        `3s3 u\�s3z3 Pz3�3 u\��3�3 P�34 u\��9�9 u\�        �34 0��9�9 0�        �3�3 u\��3�3 P�34 u\��9�9 u\�        �34 0��9�9 0�        �3�3 u\��3�3 P�34 u\��9�9 u\�        �34 	���9�9 	��        �34 S�9�9 S        �3�3 u\��34 P44 u\��9�9 u\�        �34 0��9�9 0�        �34 F���9�9 F��        �34 S�9�9 S        �3�3 u\��34 P44 u\��9�9 u\�        44 uT#4"4 P"4#4 t #4'4 t        4"4 u\�"4'4 P'4B4 u\�B4G4 PG4K4 u\�~7�7 u\�        K4�5 ���6[7 ���8�8 ���9�9 ���9: ��        K4�4 u#O7S7 PS7[7 u#        r4u4 u`�u4�5 W�6O7 W�8�8 W�9�9 W�9: W        �4�4 w         �4�4 0��4�4 s u #��4�4 s u #��4M5 s u #��6O7 s u #��8�8 s u #��9�9 s u #�        �4�4	 s �H$H&��6�6	 s �H$H&��67	 s �H$H&�77 p H$H&�707	 s �H$H&�0767 p H$H&�97G7	 s �H$H&��9�9	 s �H$H&�        77 u�        77 u`�        97C7 u\�C7L7 PL7O7 u\�        97O7 u`�        �9�9 u`�        
5�5 u`��8�8 u`��9�9 u`��9�9 u`�        #5A5 u�        #505 u@r �05:5 P        #5A5 0�        #5A5 u`�        A5�5 u@�9�9 u@�9�9 S        A5W5 P        A5f5
 uH�uO��f5�5
 uH�uO���9�9
 uH�uO���9�9 uH��        A5�5 �B�  �9�9 �B�          G5f5 u@�9�9 S        G5W5 P        G5f5 uH�9�9 uH        f5�5 u`��9�9 u`�        i5�5 u[��9�9 u[�        i5t5 P�9�9 P        t5�5 u\�        z5�5 u`�        z5�5 P        �9: u`�        �9: u[�:: R:: u[�        �9: P        :*: u\�        :: u`�: : R :*: u`�        : : P        �5�5 0�        �5�5 u#        �5 6 u         `:l: �o:r: P�u�        �:�: P�:6; u@�=6> u@�@�A u@BB u@JB~B u@        �:6; W�=> W>> w�>&> W&>6> R6>�> u��?�@ u�        �:�: V�: ; uT#>> q$> > uT#$        
>> q(> > uT#(        6;t< V�<�< V0=Z= Ra=�= u@o?�? V�@�@ R�A�A R�A�A u@�A�A S�AB VBB V        �:P; u�=�> u�?�@ u�@�A uBB uJByB uyB~B uDl�        �:�: uD�=
> uD�@�A uDBB uDJB~B uD        �:�: P�:�: W�@�A WBB WJB~B W        �:�: u#l#�@A u#l#        �@�A 0��A�A SBB 0�BB SJBSB 0�[BnB S        A�A 0�BB 0�[BnB 0�        A�A SBB S[BnB S        �:P; u �=�> u �?�@ u         �:6; S�=�= S>3> S3>�> W�?D@ WN@�@ W        �:; W;4; P�=�= P>&> W&>6> R6>�> u��?�@ u�        �:�= 8��=�= 8�>�@ 8��AB 8�BJB 8�        �:6; u@�=�= u@>6> u@         >&> W&>6> R6>�> S�?I@ SN@�@ S        6>P> s P>�> uT�>�> u@�#0��?G@ uTG@N@ u@�#0�N@�@ uT        6>�> 8��?�@ 8�        6>P> 0�P>�> V�>�> P�>�> V�?%@ V%@>@ P>@A@ VN@�@ V        6>P> 0�S>�> Q�>�> u��>�> Q�?@ Q@%@ u�%@]@ Q]@p@ u�p@}@ Q}@�@ u��@�@ Q�@�@ u��@�@ Q�@�@ u��@�@ Q�@�@ u�        6>P> 1�_>�> P�?�? P�?�? 1q �$��?�? P�?�? 1q �$��?@ PN@]@ Pp@}@ P�@�@ P�@�@ P�@�@ P        �>�> P�?�? P�?�? P@%@ Pi@p@ P�@�@ P�@�@ P�@�@ P�@�@ P        g;x; Rx;�; S�;�< u@o?{? u@{?�? S�?�? u@BB u@        �<�< P�<�< Q�<a= u@�>o? u@�@�@ u@�A�A u@        �<�< R�<�= u��>o? u��@�@ u��A�A u�        >;O; u\�O;T; PT;�; u\��;�; P�;�; u\��;�; P�;�= u\��>�? u\��@�@ u\��AB u\�BJB u\�        K;O; u\O;P; p �<�< w         >;O; u\�O;T; PT;�; u\��;�; P�;�; u\��;�; P�;�< u\��<�< u`��<�= W�>o? Wo?�? u\��@�@ W�A�A W�AB u\�BB u\�B,B W        �;< S        �;0< 0�BB 0�        �;�; s 1$��;�; P�;�; t �;�; t�;�; t�;�; t�;�; s 1$��;0< u@1$�BB u@1$�        �;�; u\��;�; P�;�; u\��;�; P�;0< u\�BB u\�        �;0< 0�BB 0�        �;�; u\��;�; P�;0< u\�BB u\�        �;0< 0�BB 0�        �;�; u\��;< P<0< u\�BB u\�        <0< 	��BB 	��        <0< SBB S        << u\�<&< P&<0< u\�BB u\�        <0< 0�BB 0�        <0< F��BB F��        <0< SBB S        << u\�<&< P&<0< u\�BB u\�        4<?< uT#?<B< PB<C< t C<G< t        4<B< u\�B<G< PG<b< u\�b<g< Pg<k< u\��?�? u\�        k<�= ���>{? ���@�@ ���A�A ��B,B ��        k<�< u#o?s? Ps?{? u#        �<�< u`��<�= W�>o? W�@�@ W�A�A WB,B W        �<�< w         �<�< 0��<�< s u #��<= s u #�=m= s u #��>o? s u #��@�@ s u #��A�A s u #�        �<�<	 s �H$H&��>?	 s �H$H&�?,?	 s �H$H&�,?1? p H$H&�4?P?	 s �H$H&�P?V? p H$H&�Y?g?	 s �H$H&��A�A	 s �H$H&�        &?4? u�        &?4? u`�        Y?c? u\�c?l? Pl?o? u\�        Y?o? u`�        �A�A u`�        *=�= u`��@�@ u`��A�A u`��A�A u`�        C=a= u�        C=P= u@r �P=Z= P        C=a= 0�        C=a= u`�        a=�= u@�A�A u@�A�A S        a=w= P        a=�=
 uH�uO���=�=
 uH�uO���A�A
 uH�uO���A�A uH��        a=�= �"�  �A�A �"�          g=�= u@�A�A S        g=w= P        g=�= uH�A�A uH        �=�= u`��A�A u`�        �=�= u[��A�A u[�        �=�= P�A�A P        �=�= u\�        �=�= u`�        �=�= P        B,B u`�        B'B u[�'B+B R+B,B u[�        B+B P        ,BJB u\�        2B<B u`�<B@B R@BJB u`�        2B@B P        �=�= 0�        �=�= u#        
> > u         �B�B P�B�C W�C*D W.DCD W        �B*D 
G�.DCD 
G�        �B�B P�B�B S�B*D ��.DCD ��        �B�B P�B*D �@.DCD �@        �B*D 0�.DCD 0�        �B�C S�C�C �\��CD SD&D �\�&D(D S(D*D �\�.DCD �\�        C&D �L        C&D	 ���@"�        C&D ��        C�C W�C&D W        :CNC �L        :CNC	 ���@"�        :CNC ��        :CNC W        wC�C S�C�C �\��CD SD&D �\�        zC�C �W��CD �W�DD PD&D �W�        zC�C R�CD R        �CD �W�DD PD&D �W�        �CD R        �C&D 	��        �CD r�        DD QD&D s�        .DCD �\�        4D>D �W�>DBD RBDCD �W�        4DBD P        �DE �!E.E V.E2E t SE�E ��E�E V�EF �FF VFG �        EME WMESE ���SE�E W�E�E ��E�E ����EG W        EE 0�!E2E R2ESE �\SE�E 0��E�E 1��EF 0�FF 2�FG 0�        EE PEE qSEfE qfEgE � #�E�E q        uEE PE�E QF,F P,FIF �\�FG �\        SEfE QfE�E � �EG �         uE�E -��EG -�        �E�E -�FG -�        F,F P,FIF �\�FG �\        �E�E X��F�F X�        �E�E Q�F�F �\        �E�E +��EF +�UF�F +�        �E�E QUFnF QnF�F �\        �E�E 0��EF 0��F�F 0�        �E�E Q�F�F Q�F�F �\        �E�E x��EF x��F�F x�        �E�E Q�F�F �\        !ESE �X        !EME WMESE ���        !E.E V.E2E t         3E=E s �\�=EKE SKERE �RESE ��\�        3E?E u �\"�?ENE UNERE �RESE ��\"�        �E�E S�E�E �D�E�E �        �E�E U�E�E �        �E�E V        �E�E �X        �E�E W�E�E ��E�E ���        PGnG � nG�G U�G�G � �G�G U        PGnG �nG�G Q�G�G R�G�G Q�G�G P�G�G Q�G�G P�G�G Q        PG�G ��G�G V�G�G ��G�G V        eGnG � nG�G S�G�G U�G�G S�G�G U�G�G S        �G�G
 �
 @0.��G�G p 0.��G�G
 �
 @0.�        �G�G 
 @�        �G�G �         HH �HH P���'I1I Q�W�        @HPH �H        SH4J D��J�J D�        VH�H V�H�H t	���H�H P�H�H t �H�H t�H�H t�H�H t�HI tII tI1I PZIjI p�jI�I P�I�I t�I�I t�I�I t�I�I t�I�I t�I�I V�I�I P�I�I p~��IJ PJ*J p�*J4J P�J�J p��J�J P        qH�H R�H�H ��tI�I ��        �H�H P�H�H t �H�H t�H�H ������0+�+( �tI�I ������0+�+( �        H�H �#l�tI�I �#l�4J�J �#l��JK �#l�        'H*H P*HMH V4J�J V�JK V        'H@H �#l#4JIJ P        4J�J 0��J�J W�J�J W�J�J 0��J�J W�J�J 0�        QJ�J 0��J�J 0��J�J 0�        QJ�J W�J�J W�J�J W        VH4J J��J�J J�        VH�H Q�H�H �@tI�I �@        �I�I V�I�I v~�        �I�I	 q 
 @0.�        �HI V        IZI 0�        II �#         ITI S         I1I P        I I �L�� I,I	 �L�R��,I?I	 �L�V��?IUI	 �L�V��UIZI
 �L�p��         IZI ��          $I?I S        $I1I P        $I?I �L        H�H �tI�I �4J�J ��JK �        KnK �        /KIK vIK�K �L�K�K P�K�M �L        9KHK w ��HKgK W        �K�K W�K�L �H�L�L W�L$M �H�M�M �H        �K�K R�K�L �D�L�L R�L�L �T�L$M �D�M�M �D        �KeL v� ��L�M v� ��M�M �#l��M�M v� ��M�M �#l�        �K�K P�K�K Q�K�K �H�L�L �H$M9M Q9M�M �H�M�M �H        �K�K v� #$M5M v� #        $M�M 0��M�M R�M�M �@�M�M �@�M�M 0��M�M �@�M�M 0�        DM�M 0��M�M 0��M�M 0�        DM�M R�M�M �@�M�M �@�M�M �@        �KL W�L$M W�M�M W        �K�K Q�K'L �P'L,L t	��,L/L t	��/L0L t	��0L1L t	��1L7L t	��7LGL t	��GLKL t	��KLNL t	��NLOL t	��OLXL t	��XL^L t	���L$M �P        �K�K �P�K�K P        �KL W�L$M W�M�M W        L�L ���L$M ���M�M ��        L�L �L�L$M �L�M�M �L        �KeL V�L$M V�M�M V        �K�L 0��L$M 0��M�M 0�        �KL v        'L^L W        'L3L Q        'LBL	 S��T��BL^L S��        'L^L �~�          )L^L W        )L3L Q        )L^L S        BLQL RQL^L �P        BL^L �H        BL^L ��          BL^L S        �L�L R�LM �TM$M �D        �L$M �H        �L�L	 S��T���L$M S��        �L$M ��          �L�L R�LM �TM$M �D        �L$M �H        �L$M S        M$M W        MM QM$M �P        M$M �/�          M$M S        �L�L R�L�L �T        �L�L �H        �L�L	 S��T���L�L S��        �L�L ��          �L�L R�L�L �T        �L�L �H        �L�L S        �L�L V        �L�L 0�        �L�L v        �KeL V�L�M V�M�M ��M�M V�M�M �        cN�N �        cN�N �        cNzN QzN�N �        cNzN PzN�N �        �N�N ��N�N P����O�O W�P��O�O W�P�        OO POQO VQO�P ��Q Q ��        O�P D�Q Q D�        OHO QHOYO �@YO�O Q�O�O Q�O*P Q:P@P P@PaP QaPuP q~�uP�P QQQ q�Q Q Q        :OHO RHO�P �KQ Q �K        :OmO ��O P �        �NmO �#l��O
P �#l��PQ �#l� QXQ �#l�        �N�N P�NO W�PQ W QXQ W        �N O �#l#�P�P P        �P�P 0��P�P P�PQ S Q"Q S"Q$Q 0�$Q5Q S=QHQ 0�        �PQ 0� Q"Q 0�$Q5Q 0�        �P�P P�PQ S Q"Q S$Q5Q S        O�P J�Q Q J�        OmO W�OiP WQ Q W        PP PP*P p~�*P@P �@2�        aPiP	 w 
 @0.�        �O�O S        �O�O 0�        �O�O �#        �O�O V        �O�O Q        �O�O �L���O�O	 �L�P���O�O	 �L�S���O�O	 �L�S���O�O
 �L�p��        �O�O �D�          �O�O V        �O�O Q        �O�O �L        �NmO ��O
P ��PQ � QXQ �        �Q�Q ��QR V�W�        �QR URR �#        �Q�Q u ����Q�Q P�QR u ���RR �#���        �Q
R S
RR �        �QR URR �#        3RXR �        3RXR �        3RJR QJRXR �        3RJR PJRXR �        �R�R ��R�R �X�R�R P�R�
S/S �/SOS �XSS]S V�W�]SaS �aS�S �X�S�S P�R�        �R�R � �RS S
S/S � /S]S S]SaS � aS�S S        S#S
 �
 @0.�#S(S p 0.�(S]S
 �
 @0.�        S]S 
 @�        S]S �        �S�S ��S�S P���UU V�V�U U W�V�        	TT PTV ���V�V ��        TV (��V�V (�        TuT SuT�T t	���T�T P�T�T t �T�T t�T�T t�T�T t�T�T t�T�T t�TU P%U:U p�:UpU PpUqU tqUtU ttUwU twUzU tzU~U t�U�U S�U�U P�U�U p~��U�U P�U�U p��UV P�V�V p��V�V P        T,T �G        WTjT P�R�        �S�T �#l�DUaU �#l�V�V �#l��V�V �#l�        �S�S P�S{T WV�V W�V�V W        �S�S �#l#VV P        VkV 0�kV�V V�V�V V�V�V 0��V�V V�V�V 0�        !V�V 0��V�V 0��V�V 0�        !V�V V�V�V V�V�V V        TV J��V�V J�        TT PTbT �#bTV ���V�V ��        eUhU ShU�U s~�        �U�U ��
 @0.�        �T�T S        �T%U 0�        �T�T �#        �TU W        �TU P        �TU	 �@�S��UU	 �@�S��U%U
 �@�p��        �T%U ��          �TU W        �TU P        �TU �@        �S�T �DUaU �V�V ��V�V �        MWjW V�W�        MWoW �        MW_W Q_WoW �        MW_W P_WoW �        �W�W ��W�W P����X�X W�P��X�X W�P�        �W0X V0XrY ���YZ ��        �WrY (��YZ (�        �W'X Q'X8X ��8X~X Q�X�X Q�X
Y QYY PYGY QGY\Y q~�\YrY Q�YZ q�ZZ Q        X'X R'XLX W�X Y W Y0Y P0Y5Y W        XrY �@�YZ �@        �WLX �#l��X�X �#l�rY�Y �#l�ZHZ �#l�        �W�W P�WX WrY�Y WZHZ W        �W�W �#l#rY�Y P        rY�Y 0��Y�Y SZZ SZZ 0�Z%Z S-Z8Z 0�        �Y�Y 0�ZZ 0�Z%Z 0�        �Y�Y SZZ SZ%Z S        �WrY J��YZ J�        �W�W P�WX �#XrY �L�YZ �L        �X�X P�X
Y p~�
Y Y ��2�        GYrY
 �L
 @0.�        mX�X S        �X�X 0�        �X�X �#        �X�X V        �X�X Q        �X�X �H���X�X	 �H�P���X�X	 �H�S���X�X	 �H�S���X�X
 �H�p��        �X�X ��          �X�X V        �X�X Q        �X�X �H        �WLX ��X�X �rY�Y �ZHZ �        �Z�Z V�W�        �Z�Z �        �Z�Z Q�Z�Z �        �Z�Z P�Z�Z �        [[ P[/[ W1[�[ W�[(\ W        [-[ s #-[0[ u#0[1[ t#1[E[ s #        1[�[ 0��[�[ P�[�[ ud�[�[ �\�[�[ 0��[�[ ud�[�[ 0�\\ ud        L[�[ 0��[�[ 0�\\ 0�        L[�[ P�[�[ ud�[�[ �\�[�[ ud\\ ud        H\J\ PJ\_\ Wa\] W]X] W        H\]\ s #]\`\ u#`\a\ t#a\u\ s #        a\�\ 0��\] P]] ud]] �\]] 0�]!] ud!]*] 0�2]H] ud        |\] 0�]!] 0�2]H] 0�        |\] P]] ud]] �\]!] ud2]H] ud        x]z] Pz]�] W�]^ W^S^ W        x]�] s #�]�] u#�]�] t#�]�] s #        �]�] 0��]�] P�]^ ud^^ �\^^ 0�^^ ud^%^ 0�-^C^ ud        �]^ 0�^^ 0�-^C^ 0�        �]�] P�]^ ud^^ �\^^ ud-^C^ ud        `^q^ �}^�^ P����_�_ W�P�
`` W�P�        �^�^ P�^�_ ��`;a ��        �^_ S        �^�^ w40.�        �^�^ P�^�^ pb��^�^ sv w�4H$0)( �        �^�_ V`�` V�`a V a;a V        _Q_ P�`�` P�`�` �� a/a P        +_/_ Q/_�_ ���_` ��`�` ���`�` ���`;a ��        l_�_ 0��_�_ P`X` 0�        t^�_ W`;a W        +_/_ Q/_;a ��        +_a_ v s "��`�` v s "� a;a v s "�        +_�_ V`�` V�`a V a;a V        +_Q_ P�`�` P�`�` �� a/a P        Q_f_ ��        Q_a_ v s "�        Q_f_ V        l_�_ S`�` S�`a Saa s�a a �H#�        l_�_ V`�` V�`a V        k`n` Rn`�` ���` a ��        k`�` 0��`�` S�` a 1�        �_�_ S        �_` 0�        �_�_ w        �_�_ R�_
` ��        �_` ��        �_�_ �����_�_
 ���P���_
`
 ���S��
``
 ���S��`` ���p��        �_` ��          �_�_ R�_
` ��        �_
` ��        �_
` ��        �a�a ��a�a P���cc W�P�$c'c W�P�        �a�a P�a
c ��9c[d ��        �a-b S        �a�a w40.�        �a�a P�a�a pb��a�a s$v w�4H$0)( �        b�b V9c�c V�c#d V@d[d V        *bkb P�c�c P�cd ��@dOd P        EbIb QIb�c ���c�c ���cd ��d@d ��@d[d ��        �b�b 0��b�b P9cxc 0�        �ac W9c[d W        EbIb QIb�b ���b9c ��9c�c ���c�c ���cd ��d@d ��@d[d ��        Eb{b v s "��cd v s "�@d[d v s "�        Eb�b V9c�c V�c#d V@d[d V        Ebkb P�c�c P�cd ��@dOd P        kb�b ��        kb{b v s "�        kb�b V        �b�b S9c�c Sd&d S&d3d s�3d@d �H#�        �b�b V9c�c Vd#d V        �c�c R�c�c ��d@d ��        �c�c 0��c�c Sd@d 1�        �b�b S        �b9c 0�        �b�b w        �bc Rc$c ��        �b9c ��        �b�b �����bc
 ���P��c$c
 ���S��$c3c
 ���S��3c9c ���p��        �b9c ��          cc Rc$c ��        c$c ��        c$c ��        �d�d 	���d�d P�d�d 	���d�d P�d�d 	���d�d P�de 	��        �d�d R�d�d R        �d�d P�d�d P        �d�d P        �d�d R        �d�d P        eKe VKeLe � Le�e V�e�e � �e�e V�e�e � �e�e V        e/e 	��Le[e 	��[ebe P�e�e 	���e�e P�e�e 	��        Le[e P�e�e P        [ebe P�e�e P        Xe[e R        �e�e P        �e�e P        /eJe SJeLe �be�e S�e�e ��e�e S�e�e ��e�e S        /eLe 	��be�e 	���e�e 	���e�e 	��        /eAe 	��be{e 	��{e}e P�e�e 	���e�e P�e�e 	��        be{e P�e�e P        {e�e P�e�e s�e�e �#�e�e P        xe{e Q        �e�e P        �e�e P        ff PfGf Wpf�f W        :fGf Spf�f S�f�f �T        :fGf 0�pf�f 0��f�f S�f�f s��f�f S�f�f P�f�g �\�g�g V�g|h �\|h�h V�hi �\        :fGf 0�pf�f 0��fkg �Xngyg Pyg8h �X;h|h V|h�h �X�hi V        :fGf 1�pfi 1�        �g�g	 w 2$�";huh W|h�h	 w 2$�"�h�h	 w 2$�"�hi W        :f;f t ;f?f t?fyg ��yg�g P�g�g t �g�g t�gSh ��ShZh PZh[h t [h_h t_hi ��        :f?f P?fsf ��sf{f P{f�g ���g�g P�gZh ��Zh_h P_h�h ���h�h Q�hi ��        ~f�f P        pfsf ��sf{f P{f�g ���g�g P�gZh ��Zh_h P_h�h ���h�h Q�hi ��        ~f�f 0��f�f V        �f�f P        �f�f W        GfVf 4�        GfVf �(        GfVf �(        gg Pg g W gGg SGg�g W�h�h W        �fg	 s 2$�"        g g 1� g�g V�h�h V         g,g v 2$w "2$�"        Gg�g ���g�g P�gh ��|h�h ��        Ng`g P�h�h P        Zg`g 1�        �h�h P        vgyg ��yg�g P�g�g t �g�g t�gh ��|h�h ��        vg�g ���g�g P�gh ��|h�h ��        �g�g R�gh R|h�h R�h�h �T�h�h R        �g�g ���gh ��|h�h ��        �g�g 	���gh 	��|h�h 	��        �g�g 	���g�g P|h�h 	���h�h P�h�h 	��        �g�g Q|h�h Q        �g�g P�h�h P        �g�g P        �h�h Q        �h�h P        hZh ��Zh_h P_h|h ���h�h ���h�h Q�hi ��        ;huh W�hi W        PhSh ��ShZh PZh[h t [h_h t_hgh ���hi ��        PhZh ��Zh_h P_hgh ���h�h ���h�h Q�hi ��        �h�h ���h�h Q�hi ��        +i.i P.iqi �T�k�l �T�l�l �T�l m �T        IiLi PLiqi W�k�k W�k�l �P�l�l W�lm �P        Iiqi 0�qi�j V�j^k V�k�k V�k�k 0��k-l V-l6l v�6l�l V�l�l V�l�l 0��lm V        Iiqi 0�qi�k �T�k�l 0��l�l �T�lm 0�        Iiqi 0�qisj �\xj�k �\�kfl 0�fl�l 1��l�l �\�lm 0�        IiLi ��LiRi PRim ��        Iiai Sai�k ���k�k S�k�k t �km ��        �k�k P        �k�k S�k�k t �k�l ���lm ��        �k�k 0��kFl S�l�l 0�        ll P        l#l �T        iqi �$�k�l �$�lm �$        qi�k ���l�l ��        qi�k ���l�l ��        qi�k 	���l�l 	��        qi�i 	���i�i P�j�j 	���j�j Pk k 	�� k3k P3kDk 	��        �j�j Sk3k S        �j�j P k3k P        �j�j P        k3k S         k3k P        �i�i ���i�i ���i�i ���j�j ��  �j�j ���j�j ��  �jk ��kk �   �k�k ���k�k ��  �k�k ���k�k �           �i�i ���  �i�i ��  �i�i ���  �i�i �   �j�j ���  �j�j ��  �j�j ���  �jk �   3kDk ���  �k�k ��  �k�k �   �l�l ���          �i�j ���jk ��3k�k ���l�l ��        �i�j 	���jk 	��3k�k 	���l�l 	��        �i�i 	���j�j 	���j�j P3kDk 	���k�k 	���k�k P        �j�j R�k�k R        �j�j P�j�j ��k�k P        �j�j P        �k�k R        �k�k P        �i�i 0��i�i 0��i�i �L�i�j �L�jk 0�DkXk �L�k�k 0��l�l 0�        �i�j �KDkXk �K        �i�i ���jk ���k�k ���l�l ��        �i�i 	���jk 	���k�k 	���l�l 	��        �i�i 	���jk 	��kk P�k�k 	���k�k P�l�l 	��        �jk R�k�k R        kk P�k�k P        kk P        �k�k R        �k�k P        �i�i 0��ihj Rxj�j RDkLk R        �i�i Sj,j S,j<j
 �P2$�"xj�j S        Ojxj ��DkXk ��        Vjhj SDkPk S        bjhj 1�        DkPk S        �j�j 4�        �j�j �(        �j�j �(        Ll�l ��        �l�l S        �l�l s 2$w "2$�"        m�n ��n�n �        4m;m P;m/n S        )m1m P1m(o �        <m�m ����m�m R�m�m t �mn ��~n(o ���        <m/n S        |m/n S        On�n �  �n(o �          On�n �p  �n(o �p          On�n 	���n(o 	��        On\n 	��\nbn U�n�n 	���n�n U�no 	��o(o P        �n�n So(o S        �n�n Uo(o P        �n�n P        bnnn � �n�n � �n�n �?  �n�n � �n�n �?          \nbn �
  bnnn �5  nn|n �  �n�n �5  �no �
          \n�n �  �no �          \n�n 	���no 	��        \nnn 	���n�n 	���n�n 	���n�n P�no 	��        �n�n �        �n�n P        �n�n �        rn|n 2�        rn|n �        rn|n �        �n�n 4�        �n�n �        �n�n �        0oYq �}q�q �        Zoao Pao�p S        OoWo PWo�q �        bo�p ����p�p R�p�p t �p�p ��~�p�q ���        bo�p S        �o�p S        qYq ��  lq�q ��          qYq �  lq�q �          qYq 	��lq�q 	��        q%q 	��%q+q Ulq{q 	��{q}q U�q�q 	���q�q P        lq}q S�q�q S        {q}q U�q�q P        xq}q P        +q7q �� }q�q �� �q�q �	  �q�q �� �q�q �	          %q+q �T  +q7q �	  7qEq �U	  }q�q �	  �q�q �T          %qYq ��  }q�q ��          %qYq 	��}q�q 	��        %q7q 	��}q�q 	���q�q 	���q�q P�q�q 	��        }q�q �        �q�q P        �q�q �        ;qEq 2�        ;qEq �        ;qEq �        Yqlq 4�        Yqlq �        Yqjq �        @O �OS V���S� V�W��^� V�W�        @� ��'� �        `c P        `c p#�p#�cm p�p�mq t ��q� �@��        W� U�^� �        �� 	���� Q�� 	���� Q'�L� 	��L�^� P        �� V@�^� V        �� QL�^� P        �� P        �� � �� � �� ��  �� � �'� ��          �� ��  �� ��  �� ��  �'� ��  '�@� ��          �� �  �@� �          �� 	���@� 	��        �� 	���� 	���� 	���%� P'�@� 	��        �'� �        �%� P        �'� �        �� 2�        �� �        �� �        `�o� �o�s� V���s�� V�W��~� V�W�        `�� ��G� �        ���� P        ���� p#�p#����� p�p����� t ������ �@��        w��� U��~� �        ��ƀ 	��ƀ̀ Q�� 	���� QG�l� 	��l�~� P        �� V`�~� V        �� Ql�~� P        �� P        ̀Հ � �� � �� �  �0� � 0�G� �          ƀ̀ �[  ̀Հ �  Հ�� �Y  �G� �  G�`� �[          ƀ� �  �`� �          ƀ� 	���`� 	��        ƀՀ 	���� 	���0� 	��0�E� PG�`� 	��        �G� �        0�E� P        '�G� �        ـ�� 2�        ـ�� �        ـ�� �        ���� P���� u@���� ����ގ u@ގ� t��'� u@        ���� P���� uL���� �D��ގ uLގ� tH�'� uL        �� � V ��� u����� ����ގ u�ގ� t��� u��� V�'� u�        ��9� 0�t��� 1��� 0�        ��9� 0�c�� w ��� u�t��� w(���� u��� 0�        ā�� u����� ����ގ u�ގ� t��'� u�        �9� 0��� VǇ u�        �9� 0����� v���Ǉ 0��� 0�        �T� 1�T�^� uP���� uP��� 1��"� uP"�<� 0���C� 1�C�I� uP[�e� uPn��� 1�:�� 1���ԉ 1���&� 1�V�� 1�=��� 1����� 1�W��� 1�        �9� 0���Ǉ 1�        &�(� V(��� uH���� �@��ގ uHގ� tD�� uH        ���� u �� u         āׁ u\�ׁ� P��� u\����� �T���ގ u\�ގ� tX��'� u\�        ΁ׁ u\ׁ� p ��� p         āׁ u\�ׁ� P�� u\��� u`���� P���� u`����� �X���ގ u`�ގ� t\��� u`��� u\��	� u`�        �� u`���� P���� u`����� �X���ގ u`�ގ� t\��� u`��	� u`�        ��� p         +�9� V9�E� P���� uD#���ł P        +�9� u v "L�H$H&���ł u p "L�H$H&�        ؆� S�<� Sԉ�� S�.� S        ؆�  ��<�  �ԉ��  ��.�  �        ؆� u@�$� Q$�<� u@ԉ�� u@�.� u@        0��� uT��<� uT        3�j� Qj�v� u�v��� Q���� q����� Q��ǈ u�ǈۈ Qۈ� u��� Q�� u��+� Q+�<� u�        <�j� P���� Pǈۈ P�� P��	 w q �$��� P�+� P        v��� Pňǈ P�� P�� P7�<� P        f��� u���:� u���� u�ԉ�� u�&�V� u��=� u�        f��� u���:� u���� u�ԉ�� u�&�V� u��=� u�        f��� 	����:� 	����� 	��ԉ�� 	��&�V� 	���=� 	��        f�z� 	��z��� P���� 	������ P�!� 	��f�|� 	��|��� P        ���� Rf�x� R        ���� P|��� P        ���� P        f�x� R        z��� u����� u����� �  ��҆ u�҆Ն ��*  �!� u�0�:� �   L�f� �   &�<� u�<�V� ��*          z��� �z  ���� �   ���� �{   ���� �z  ���� �{   ��Ն ��*  �� �z  �:� �   <�f� �   &�V� ��*  .�=� �{           z��� u����� u��!� u�        z��� 	����:� 	���f� 	��ԉ�� 	��&�V� 	���=� 	��        z��� 	������ 	���0� 	��0�5� P5�:� u<�L� 	��L�a� P        !�0� R<�H� R        0�5� P5�:� uL�a� P        -�0� P        <�H� R        l��� u�        ��� u���ă u�        ��� u���ă u�        ��"� 	��:�� 	����ԉ 	������ 	��=�F� 	��        ���� 	����� P��� 	��:�O� 	��O�h� P��� 	���!� P        :�O� R��� R        O�h� P�!� P        L�O� P        ��� R        ��� u��� u�'�0� u��� u���� �#  U�h� �"  w��� u����� ��#  <�V� �#  V�l� u�l��� ��#          ��� ��!  �� ��"  �'� ��"  '�0� ��#  ă� ��!  �� ��"  �� ��"  U�]� ��!  ]�w� ��"  w��� ��#  !�V� ��"  V��� ��#          ��� u�ă� u�U�h� u�        ��"� 	��U�� 	����ԉ 	��!��� 	��=�F� 	��        ��� 	��ă�� 	����� PU�]� 	��!�<� 	��<�Q� P        ��� R!�8� R        ��� P�� u<�Q� P        ���� P        !�8� R        5�d� S���� SǇ� S=�F� S        �$� u�'�0� u�]�h� u�w��� u�V��� u�        �0� 	��]��� 	��V��� 	��        �0� 	��]��� 	������ PV�l� 	��l��� P        w��� RV�h� R        ���� Pl��� P        ���� P        V�h� R        5�ă �#  ��� �#  ��ԉ �#  =�F� �#          5�ă :���� :���ԉ :�=�F� :�        5�ă uH��� uH��ԉ uH=�F� uH        [��� W���� Q���� Q        [��� u`����� u`�        d��� S���� S        ���� ��$  ���� ��$          ���� p r "�        ���� u`����� u`�        ���� S���� S        ���� pt����� pt�        ���� S        ���� pt�        ���� p s "�        �� 0�        ��� u\��	� P	�� u\�        ��ă u���ԉ u�        ���� R��ȉ R        ���� 1�        ��ȉ R        �"� u`�        ���� P��&� uT        ���� 0���&� S        ��&� u�        ��&� u�        ��&� 	��        �� 	��&�<� 	��<�H� PH�`� 	������ 	������ P        &�8� P���� P        &�8� P        <�H� P���� P        ���� R        ˊ׊ u�Z�`� u�o�~� �<)  �&� �<)          ˊ �(  ˊ׊ �2)  ׊� �)  H�Z� �(  Z�t� �2)  t�~� �)  ��� �)  �&� �2)          ׊ u�H�`� u�        &� 	��H��� 	����&� 	��        ׊ 	��H�o� 	��o�t� P�� 	���&� P        `�o� P�� P        o�v� Pv�~� u�&� P        l�o� R        �� P        �� u���� P��� u���� u�        ��� u�        ��ŋ Pԋ� P        ��ŋ 1�        ԋ� P        �#� u�#�*� P*�+� t +�/� t/�I� u�V��� u�        �*� u�*�/� P/�I� u�V��� u�        ��Ն u�&�V� u�.�=� u�        ��Ն 	��&�V� 	��.�=� 	��        ��҆ 	��҆Ն P؆� P�"� P&�<� 	��<�V� P.�=� 	��        Æ҆ R&�8� R        ҆Ն P<�V� P        φ҆ P        &�8� R        ��� u�ԉ�� u��.� u�        ԉ� R�%� R        �� 1�        �%� R        V�Y� u�Y�a� Pa��� u�        ~��� u�        ���� u����� P���� t ���� t��، u�F��� u�        ���� u����� P��، u�F��� u�        }��� u�        �� u��� P��� t ��� t�� u�W��� u�        �� u��� P�� u�W��� u�        F�I� u�I�Q� PQ��� u�        W�Z� u�Z�b� Pb��� u�        6�<� 4�        6�<� u$        6�<� u$        <��� u����� ������ u�̎ގ u�ގ� t��� u�        <��� u����� ������ u�̎ގ u�ގ� t��� u�        b��� u`����� �X�̎ގ u`�ގ� t\��� u`�        e��� u[����� �S�̎ގ u[�ގ� tW��� u[�        e�p� P�� P        p��� u\����� �T�̎ގ u\�ގ� tX�        v��� u`����� �X�̎ގ u`�ގ� t\�        v��� P���� u\<����� �T<�̎ӎ P        ̍W� uP        ̍ٍ 1�ٍG� uTI�W� uT        ٍW� u�        ٍW� u�        �W� u�        '�W� u�        .�<� RI�Q� R        6�<� 1�        I�Q� R        e�|� u`�|��� P���� u`���̎ u`�        ���� P        ���� p 	�)�        ���� u`�        ��� 0���̎ 0�        ��ǅ u`�ǅυ Pυ� u`��� P�� u`���̎ u`�        օ� u`��� P�� u`���̎ u`�        ۅ� u`��� P�� u`�        �� -�        �� u`��� P�� u`�        �� 0�        �� pt�        �,� u\�,�V� SV��� u\����� S        /�8� P8�V� v H$H&u��H$H&u��0)( ����� v H$H&u��H$H&u��0)( �        /�V� S���� S        ���� 4�        ���� u$        ���� u$        ���� 2�        ���� u$        ���� u$        �	� u`�        ��� u[��� R�	� u[�        ��� P        �� u`��� R�'� u`�        �� P        H�I� PI�;� u@;�>� t�>��� u@���� t���ל u@        `�n� Pn�;� uL;�>� tH>��� uL���� tH��ל uL        g�Џ VЏ;� u�;�>� t�>��� u����� t����� u����� V��ל u�        g�� 0�$�X� 1����� 0�        g�� 0��/� w /�C� u�$�@� w(@�X� u����� 0�        t�;� u�;�>� t�>��� u����� t���ל u�        ��� 0�i�r� Vr�w� u�        ��� 0�I�L� v�p�w� 0���ĕ 0�        ��� 1��� uPK�U� uPg�đ 1�đґ uPґ� 0�>�� 1���� uP�� uP�;� 1��ĕ 1�A��� 1���֙ 1��͚ 1��C� 1�N�i� 1��X� 1�        ��� 0�l�w� 1�        ֏؏ V؏;� uH;�>� tD>��� uH���� tD���� uH        3��� u ���� u         t��� u\����� P��;� u\�;�>� tX�>��� u\����� tX���ל u\�        ~��� u\���� p ���� p         t��� u\����� P���� u\����� u`����� P��;� u`�;�>� t\�>��� u`����� t\����� u`����� u\����� u`�        ���� u`����� P��;� u`�;�>� t\�>��� u`����� t\����� u`����� u`�        ���� p         ۏ� V��� PK�U� uD#�g�u� P        ۏ� u v "L�H$H&�g�u� u p "L�H$H&�        ���� Sĕ� S���� S͚ޚ S        ����  �ĕ�  �����  �͚ޚ  �        ���� u@ĕԕ Qԕ� u@���� u@͚ޚ u@        ��;� uTF�� uT        �� Q�&� u�&�3� Q3�6� q�6�i� Qi�w� u�w��� Q���� u����� Q��̖ u�̖ۖ Qۖ� u�        �� PF�i� Pw��� P���� P����	 w q �$����� P̖ۖ P        &�;� Pu�w� P���� Pǖ̖ P�� P        �K� u�;�� u�ĕA� u����� u�֙� u�͚� u�        �K� u�;�� u�ĕA� u����� u�֙� u�͚� u�        �K� 	��;�� 	��ĕA� 	������ 	��֙� 	��͚� 	��        �*� 	��*�5� P;�O� 	��O�]� P��є 	���,� 	��,�A� P        ;�O� R�(� R        O�]� P,�A� P        L�O� P        �(� R        *�5� u�7�C� u�U�]� �8  n��� u����� �]C  ˔є u���� �9  ��� �9  ֙� u��� �]C          *�7� ��7  7�C� �9  C�K� ��8  U�]� ��7  ]�n� ��8  n��� �SC  ��˔ ��7  ˔� �9  �� �9  ֙� �SC  ޚ� ��8          *�5� u�U�]� u���є u�        *�K� 	��U�� 	��ĕ� 	������ 	��֙� 	��͚� 	��        *�C� 	��U�]� 	������ 	����� P�� u��� 	����� P        є�� R��� R        ��� P�� u��� P        ݔ�� P        ��� R        �C� u�        ���� u�n�t� u�        ���� u�n�t� u�        ��ґ 	���ĕ 	��A��� 	����;� 	����� 	��        ���� 	������ Pn��� 	����� 	����� P���� 	����ї P        ��� R���� R        ��� P��ї P        ���� P        ���� R        ���� u����� u�א�� u����� u����� �d;  �� �g:  '�?� u�?�G� �X<  �� �d;  �� u��;� �X<          ���� �/:  ���� �Z;  ��א �0;  א�� �N<  t��� �/:  ���� �Z;  ���� �0;  �� �/:  �'� �0;  '�G� �N<  ї� �Z;  �;� �N<          ���� u�t��� u��� u�        ��ґ 	���ĕ 	��A��� 	��ї;� 	����� 	��        ���� 	��t��� 	������ P�� 	��ї� 	���� P        ���� Rї� R        ���� P���� u�� P        ���� P        ї� R        �� SG�a� Sw�ĕ S��� S        ɐԐ u�א�� u��� u�'�G� u��;� u�        ɐ�� 	���G� 	���;� 	��        ɐ�� 	���?� 	��?�G� P�� 	���1� P        '�?� R�� R        ?�G� P�1� P        <�?� P        �� R        �t� ��;  G�ĕ ��;  A��� ��;  ��� ��;          �t� :�G�ĕ :�A��� :���� :�        �t� uHG�ĕ uHA��� uH��� uH        �I� WI�L� QA�c� Q        �L� u`�A�c� u`�        �L� SA�c� S        6�I� �Q=  A�Z� �Q=          6�>� p r "�        ;�L� u`�A�c� u`�        >�L� SA�c� S        >�L� pt�A�c� pt�        A�c� S        A�c� pt�        Z�c� p s "�        ��ĕ 0�        ���� u\����� P��ĕ u\�        L�t� u�c��� u�        S�e� Rc�x� R        _�e� 1�        c�x� R        đґ u`�        [�^� P^�֙ uT        [�^� 0�^�֙ S        ^�֙ u�        ^�֙ u�        ^�֙ 	��        ^�r� 	��֘� 	����� P��� 	��8�K� 	��K�S� P        ֘� P8�K� P        ֘� P        ��� PK�S� P        H�K� R        {��� u�
�� u��.� �A  ��֙ �A          r�{� �h@  {��� �A  ���� �iA  ��
� �h@  
�$� �A  $�.� �iA  S��� �iA  ��֙ �A          r��� u���� u�        r�֘ 	����8� 	��S�֙ 	��        r��� 	����� 	���$� P���� 	����֙ P        �� P���� P        �&� P&�.� u��֙ P        �� R        ���� P        ���� u����� P���� u�S��� u�        S��� u�        g�u� P���� P        o�u� 1�        ���� P        ͒Ӓ u�Ӓڒ Pڒے t ےߒ tߒ�� u��U� u�        ͒ڒ u�ڒߒ Pߒ�� u��U� u�        ]��� u�֙� u�ޚ� u�        ]��� 	��֙� 	��ޚ� 	��        ]��� 	������ P���� Pĕҕ P֙� 	���� Pޚ� 	��        s��� R֙� R        ���� P�� P        ��� P        ֙� R        ���� u����� u�͚ޚ u�        ���� R͚՚ R        ���� 1�        ͚՚ R        �	� u�	�� P�U� u�        .�U� u�        U�X� u�X�_� P_�`� t `�d� td��� u���C� u�        U�_� u�_�d� Pd��� u���C� u�        -�X� u�        ���� u����� P���� t ���� t��͚ u��X� u�        ���� u����� P��͚ u��X� u�        ���� u���� P�C� u�        �
� u�
�� P�X� u�        �� 4�        �� u$        �� u$        �;� u�;�>� t�C�N� u�|��� u����� t����� u�        �;� u�;�>� t�C�N� u�|��� u����� t����� u�        �;� u`�;�>� t\�|��� u`����� t\����� u`�        �;� u[�;�>� tW�|��� u[����� tW����� u[�        � � P���� P         �;� u\�;�>� tX�|��� u\����� tX�        &�;� u`�;�>� t\�|��� u`����� t\�        &�4� P4�;� u\<�;�>� tX<�|��� P        |�� uP        |��� 1����� uT��� uT        ��� u�        ��� u�        ��� u�        כ� u�        ޛ� R��� R        �� 1�        ��� R        �,� u`�,�8� P8�;� u`�c�|� u`�        <�H� P        <�H� p 	�)�        E�N� u`�        f� 0�n�|� 0�        f�w� u`�w�� P��� u`����� P�� u`�n�|� u`�        ���� u`����� P���� u`�n�|� u`�        ���� u`����� P���� u`�        �� -�        ���� u`����� P�� u`�        �� 0�        �� pt�        ܓ u\�ܓ� S�;� u\�c�n� S        ߓ� P�� v H$H&u��H$H&u��0)( �c�n� v H$H&u��H$H&u��0)( �        ߓ� Sc�n� S        c�n� 4�        c�n� u$        c�i� u$        C�N� 2�        C�N� u$        C�I� u$        ���� u`�        ���� u[����� R���� u[�        ���� P        ��ɜ u`�ɜ͜ R͜ל u`�        ��͜ P        ��� ���� V�u���b� V�W�g��� V�W���̝ V�W�        �� u`��� Q�d� u`�d�g� t\�g�̝ u`�         �� u`�� q g��� u`        L�d� u`�d�g� t\����� u`�        R�a� Sa�d� ud�d�g� t`����� S        R�Z� R���� R        ���� ud�        ���� R        ���� 	��        ���� r�        ���� V        ���� ud��� R̝ ud�        �� P        Н)� �)�`� u`��� ���V� u        ��� P��[� V`�v� V        2�6� S��� S6�F� S        ӝ6� u$`��� u$        ��� ud���� R�]� ud�]�`� t`�`�v� ud�        ���� ud��� r `��� ud        &�]� ud�]�`� t`���V� ud�        M�]� ud�]�`� t`��6� ud�        M�]� uc�]�`� t_��6� uc�        M�S� R�-� R        �$� uc�$�-� P-�6� uc�        �-� R        �6� 	��        �-� r�        �-� Q-�6� s�        ��� S6�F� S        ���� u,        ��� 0�6�V� 0�        Ğ� ud�6�V� ud�        ʞ� W6�D� WD�G� t G�H� tH�I� tI�J� t        ʞΞ p s "�Ξ֞ uds "�֞�� uLs "���� uds "��� uLs "�6�F� uLs "�        ʞΞ PΞ֞ ud֞�� uL��� ud�� uL6�V� uL        ʞ� V6�V� V        ��� W        ��� uLs "�        ��� uL        ��� V        ^�h� uc�h�l� Rl�v� uc�        ^�l� P        ���� P��Ԡ V٠&� V+�u� V        ���� p� ���Ԡ v� �٠&� v� �+�u� v� �        ���� 0���"� S٠M� Su��� P���� S��� P�
� S)�Y� S��� S�o� Sף$� S~��� Sl�z� Pz��� S���� P��ͥ S!�S� S��¦ P¦˦ S˦� P��� S��� 0��*� S*�i� Pԧ٧ S��u� Su��� P���� Sب�� P~��� P��ɩ P+�U� S        ���� P��˟ 1�� � uO ��� 0�٠� 0��� uO�d� 0�~�� 0���� P�*� uO*�ԧ 0�ԧ٧ 1�٧�� 0����� uO��� 0�+�K� 0�K�U� uO        ��˟ 0���� W٠�� W��
� Q
�j� Wj�o� 1�o�d� W~�� W�� P�˦ W˦� Q*�3� 0�3�f� Qf�٧ 1�٧� W���� W��� 1���� Q�~� 1�~��� Q���� 1���� W+�K� W        ��˟ 0�y��� uP� � uPj�z� uPף� uP$�,� uPƦ˦ uP˦� uT*�3� 0�3�m� uTԧ٧ P���� uP�� uT~��� uT        ˟ � 0� �-� uOy��� uO٠�� uO��T� uO��� uO�� 0�� � uOo�z� uOף� uO$�,� uO!�S� uOƦ˦ uOզ�� 0����� 0��� uO        ˟ � 0� �-� uTy��� uT٠� uT��� 1����� uT���� uT��)� 1�)�Y� uT��� 1��� 0�� � uTo�z� uTף� uT$�,� uT �ͥ 1�!�S� 1���Ʀ 1�Ʀ˦ uTզ�� 0����� 0���� 1�        ߟԠ v� �٠˦ v� �٧�� v� ����� v� ���&� v� �+�K� v� �        ���� u ��*� u ��U� u K�U� u         ���� u����� P���� t ���� t��֠ u�֠٠ t�٠(� u�(�+� t�+�u� u�        ���� u����� P��֠ u�֠٠ t�٠(� u�(�+� t�+�u� u�        �*� Q��0� QK�U� Q        ˦� u���� u��� P�٧ u����� u����� u�K�U� u�        (�0� P        (�U� u(        1��� u�        N�Q� u�Q�X� PX�Y� t Y�]� t]��� u�        N�X� u�X�]� P]�l� u�l�t� Pt��� u�        i�l� u�l�t� Pt��� u�        ���� u�F�V� u�        ���� u�F�V� u�        ���� u��%� u�        ��٧ 	����� 	���%� 	������ 	��        ���� 	������ 	����Ĩ P�%� 	������ 	������ P        ���� R���� R        ��Ĩ PĨ̨ u���� P        ���� P        ���� R        ���� P        ���� 	��F�~� 	��        ���� 	������ P�%� 	��F�i� 	��i�~� P        ���� PJ�h� P        ���� Pi�~� P        ���� R        V�h� P        i�~� P        ���� �X  ���� u����� u���̨ �#W  ���� u����� �#W          ���� ��W  ���� �W  ���� ��V  ��Ĩ �W  Ĩ� ��V  �%� ��W  ���� �W          ˟ߟ ud�զ� ud��� P��� ud�        ٟߟ udܦ� ud         �"� S٠M� S)�Y� S��� S!�S� S         �y� :�٠� :�!�S� :����� :��� :�         �y� v� �٠� v� �!�S� v� ����� v� ��� v� �         �� u٠� u)�H� u         �� 	���"�
 s H$H&0�٠�� 	����Y� 	����� 	��!�S� 	���� 	��        �"� S        �� u(�� t         ���� e���)� e���� e�!�S� e��� e�        ��� u(�
� t         ��� u���)� u���� u�!�S� u��� u�        �2� P!�8� P        %�2� 1�        !�8� P        2�M� u���ܢ u�F�S� u�        2�M� u���ܢ u�F�S� u�        2�M� 	����ܢ 	��F�S� 	��        2�A� 	��A�M� P��̢ 	��̢ܢ Pܢ� 	��F�S� 	��        2�A� P��Ȣ P        A�M� P̢ܢ P        >�A� R        ��Ȣ P        G�M� �[  M�Y� u�
�� u��)� ��[  ��� u���� ��[          G�M� ��Z  M�Y� ��[  Y��� ��[  ��
� ��[  
�)� ��[  ܢ� ��Z  �� ��[          G�M� u�ܢ� u�        G��� 	����)� 	��ܢ� 	���� 	��        G�Y� 	��
�� 	���$� P$�)� uܢ� 	����� 	����� P        
�� R��� R        �$� P$�)� u��� P        �� P        ��� R        u��� v� �H$p H$)����� v� �H$s H$)���� v� �H$p H$)��
� v� �H$s H$)�        a�d� u�d�l� Pl��� u���
� u�        ���� P        ���� u(���� t         @�Y� .�        @�H� u(H�L� t         "�-� u����� u�        -�R� PY�h� P        9�R� 1�        Y�h� P        F�R� u�v��� u�        F�R� u�v��� u�        F�q� 	��v��� 	��        F�U� 	��U�g� Pg�q� u��̡ 	��v��� 	������ P        F�U� P~��� P        U�g� Pg�q� u���� P        R�U� R        ���� P        [�e� �^  e�q� u�ơ̡ u�ۡ� �y_  ���� �y_          [�e� �H^  e�q� �o_  q�y� �E_  ��ơ �H^  ơ� �o_  ��� �E_  ���� �o_          [�q� u���̡ u�        [�y� 	������ 	������ 	��        [�q� 	����ۡ 	��ۡ� P���� 	������ P        ̡ۡ R���� R        ۡ� P�� u���� P        ءۡ P        ���� R        �� u��� P��� u�        2�o� �T  Ǥͥ �T  ��˦ �T  ��� �T          2�o� :�Ǥͥ :���˦ :���� :�        2�o� v� �Ǥͥ v� ���˦ v� ���� v� �        N�Q�
 p uH�#0�        N�^� u(^�b� t         ��� uP        ��� ud��	� P	�� ud�        �ͥ e���˦ e���� e�        �� u(�� t          �ͥ u���˦ u���� u�        $�6� Pɩة P        0�6� 1�        ɩة P        =�@� u�@�G� PG�H� t H�L� tL�ͥ u���˦ u���ɩ u�        =�G� u�G�L� PL�[� u�[�c� Pc�ͥ u���˦ u���ɩ u�        o��� Q��˦ Q��ɩ Q        X�[� u�[�c� Pc�ͥ u���˦ u���ɩ u�        ���� P        ���� u(���� t         ���� ud����� P��Ǥ ud�        ���� uP        ���� ud����� P���� ud�        ��Ǥ .�        ���� u(���� t         �� P�� t �� t�$� uP        �� ud��� P�,� ud�        +�:� u(:�>� t         o�z� u�$�,� u�        z��� Pͥإ P        ���� 1�        ͥإ P        ���� u���� u�        ���� u���� u�        ���� 	���!� 	��        ���� 	������ P���� u,�K� 	���� 	���!� P        ���� P�� P        ���� P���� u�!� P        ���� R        ��� P        ���� ��d  ���� u�E�K� u�Z�d� ��e  l��� ��e          ���� �d  ���� �e  ��� �e  ,�E� �d  E�d� �e  S��� �e          ���� u�,�K� u�        ��� 	��,�d� 	��S��� 	��        ���� 	��,�Z� 	��Z�_� P_�d� uS�l� 	��l��� P        K�Z� RS�h� R        Z�_� P_�d� ul��� P        W�Z� P        S�h� R        £ţ u�ţͣ Pͣ� u�        y��� ud����� W٧� ud���� P���� ud�        ��֠ ud�֠٠ t`��(� ud�(�+� t`�        ��֠ uc�֠٠ t_��(� uc�(�+� t_�        ��Ϡ PϠӠ st��� P�%� st�        f�u� u��� u�        u��� P%�8� P        ���� 1�        %�8� P        ���� uP        ���� ud����� P���� W        ̨Ϩ u�Ϩר Pר� u�        �� 0�        ��� u(���� t         ]�g� uc�g�k� Rk�u� uc�        ]�k� P        ��˪ �˪�� u�z� u��� u        ���� ���� u        ��֪ V֪<� u`�<�?� t\�?�� u`�        ���� v         �˫ �wi          �˫ �fi          �˫ 	��        ��� 	��?�K� 	��K�P� P\�n� 	��n�z� Pz��� 	��        ?�K� PK�P� u\�b� Pb�z� u        K�P� Pn�z� P        H�K� R        \�b� Pb�z� u        �
� �wi P�X� �wi X�\� ��k  ���� �wi ��˫ ��k          ��� �j  �
� �k  
�� �k  P�\� �k  z��� �j  ��˫ �k          ��?� �wi  P�\� �wi  z�˫ �wi          ��?� 	��P�\� 	��z�˫ 	��        ��
� 	��P�X� 	��z��� 	������ 	����ƫ P        P�X� u���� u        ��ƫ P        ���� u        �� 2�        �� u$        �� u$        '�<� u`�<�?� t\����� u`�        *�<� ud�<�?� t`����� ud�        *�2� R���� R        ���� ud�        ���� R        ���� 	��        ���� r�        ���� Q���� s�        ӫݫ ud�ݫ� R�� ud�        ӫ� P        �;� �;�l� ur�� u��[� u        �� ��[� u        �F� VF��� u`����� t\���[� u`�        �� v         X�;� �xn          X�;� �gn          X�;� 	��        X�l� 	������ 	������ P̬ެ 	��ެ� P��� 	��        ���� P���� u̬Ҭ PҬ� u        ���� Pެ� P        ���� R        ̬Ҭ PҬ� u        r�z� �xn ��Ȭ �xn Ȭ̬ ��p  �,� �xn ,�;� ��p          l�r� �o  r�z� �p  z��� �p  ��̬ �p  ��� �o  �;� �p          l��� �xn  ��̬ �xn  �;� �xn          l��� 	����̬ 	���;� 	��        l�z� 	����Ȭ 	����� 	���,� 	��,�6� P        ��Ȭ u�&� u        ,�6� P        �&� u        ���� 2�        ���� u$        ���� u$        ���� u`����� t\���� u`�        ���� ud����� t`���� ud�        ���� R��� R        ��� ud�        ��� R        ��� 	��        ��� r�        �� Q�� s�        C�M� ud�M�Q� RQ�[� ud�        C�Q� P        `��� ���ܭ u�Z� uh�ˮ u        `��� ���ˮ u        v��� V��� u`��� t\��ˮ u`�        v�}� v         ȭ�� �ys          ȭ�� �hs          ȭ�� 	��        ȭܭ 	���+� 	��+�0� P<�N� 	��N�Z� PZ�h� 	��        �+� P+�0� u<�B� PB�Z� u        +�0� PN�Z� P        (�+� R        <�B� PB�Z� u        �� �ys 0�8� �ys 8�<� ��u  ���� �ys ���� ��u          ܭ� �t  �� �u  ��� �u  0�<� �u  Z�h� �t  ���� �u          ܭ� �ys  0�<� �ys  Z��� �ys          ܭ� 	��0�<� 	��Z��� 	��        ܭ� 	��0�8� 	��Z�h� 	������ 	������ P        0�8� u���� u        ���� P        ���� u        ��� 2�        ��� u$        ��� u$        �� u`��� t\�h��� u`�        
�� ud��� t`�h��� ud�        
�� Rh��� R        h��� ud�        h��� R        h��� 	��        h��� r�        s��� Q���� s�        ���� ud����� R��ˮ ud�        ���� P        �	� P	��� uP��� uP��h� uPq��� uP��� uP0�L� uP[�^� uPg�~� uP        �	� p� �	��� uP#J���� uP#J���h� uP#J�q��� uP#J���� uP#J�0�L� uP#J�[�^� uP#J�g�~� uP#J�        �G� 0�G�r� Pr��� Sn�u� P�� 	��/�2� P��̴ P̴մ Sմ� P�� S���� S���� P���� S̶ٶ Pٶ� S0�;� 0�;�=� P=�B� S[�g� S        ���� w @)���� w @)����� w @)���� w @)�0�E� w @)�[�~� w @)�        �ʯ uH��� uH��� uH0�Q� uH[�y� uH        ,�5� P5��� uO���� 1��� uO��� 0����� 1���� uO�� tK��� uO���� 0���� uO�u� 0����� uO��h� 0�h�q� 1�q�� 0��-� uO-�0� tK0�;� P;�B� uOB�~� 0�        ,�J� 0�N��� uL��� uL��� uL0�;� 0�;�Q� uL[�~� uL        ���� 0���ʯ uN��ʵ 0�ʵ#� uN*��� uN���� 1����� uN��� uNB�I� uN[�g� uNg�~� 1�        ���� 0���ʯ uD�Z� uD��� uD�� t@��� uD�� � uD�� uDu��� uD2��� uD���� uD��� uD)�U� uD�� uD��ʵ 0�ʵ� uD*��� uD��-� uD-�0� t@B�g� uD        ʯ� uT�� tP��� uT��� uT�-� uT-�0� tPQ�[� uT~��� uT        ٯ�� 0���� S��� S���� 0��� S�u� 0�Q�[� 0�        ٯ� 0��ʰ W�s� Ws��� Q���� 0����� W�� Q�u� WQ�[� W        �� P�� u��� t���� u��u� u��-� u�-�0� t�Q�[� u�        �� P�� u@�� t���� u@�u� u@�-� u@-�0� t�Q�[� u@        �� 0��ٰ V��� V���� 0����� V��� V���� V�� V�� r ��u� VQ�[� V        �� 0����� 0�m��� P��� P        ��� W�� u��� uP#N��� tL#N���� uP#N����� W���� u���� uP#N���� u��F� uP#N�F�u� u��-� uP#N�-�0� tL#N�Q�[� u�        ܮG� SG��� u ��� u 0�2� S2�B� u         ��� W��#� s        �� u��	� V	�� u��� t���� u����� V���� u���� V�u� u�u�� V�-� u�-�0� t�0�Q� VQ�[� u�[�~� V~��� u�        �� u��#� P#�5� u�5�=� P=�� u��� t��-� u�-�0� t�0��� u�        2�5� u�5�=� P=��� u���� u���� u�;�Q� u�[�~� u�        o��� u����� u�        ���� u����� u�        ���� u����� P���� u����� u�        ʯ� ud��� t`���� ud���� ud��-� ud�-�0� t`�Q�[� ud�~��� ud�        ӯٯ udu��� ud        n�u� P�� 	��        ��� uT��� uT�F� uT        ��� uP#N���� uP#N��F� uP#N�        �� u��� uu��� u        �A� 	��A��� S��� 	���#� Su��� 	����� S        ��� uu��� u        ��� uP#N�u��� uP#N�        ��� uTu��� uT        A��� S�#� S��� S        R�Z� u��� u�        Z�� P���� P        f�� 1�        ���� P        s�� u����� u�        s�� u����� u�        s��� 	����� 	��        s��� 	������ P���� u�)� 	����̲ 	��̲� P        s��� P��Ȳ P        ���� P���� u̲� P        ��� R        ��Ȳ P        ���� �}  ���� u�#�)� u�8�E� �~  S�k� u�k�u� �؂  ��� u���� �؂  ,�F� �~          ���� �Q}  ���� �x~  ���� �N~  �#� �Q}  #�=� �x~  =�S� �N~  S�u� �΂  �� �΂  �F� �x~          ���� u��)� u�        ���� 	���u� 	���� 	���F� 	��        ���� 	���8� 	��8�=� P�,� 	��,�A� P        )�8� R�(� R        8�=� P=�E� u,�A� P        5�8� P        �(� R        �#� u�#�+� P+�2� u�        P��� �.y  ��� �.y          P��� uT��� uT        P��� u���� u�        ;�E� PE�F� t F�J� tJ�U� uD        ;�E� ud�E�J� PJ�Z� ud�        ���� u����� u�        ���� RZ�h� R        ���� 1�        Z�h� R        ���� u�v��� u�        ���� u�v��� u�        ��س 	��v��� 	��        ���� 	����ҳ Pҳس u��� 	��v��� 	������ P        ���� Rz��� R        ��ҳ Pҳس u���� P        ���� P        ���� R        Ƴг ��  гس u��� u�"�)� �	�  \�u� �	�          �2� �Ձ  Ƴг �؀  гس ���  س� �Ձ  ��� �؀  �)� ���  F�u� ���          Ƴس u���� u�        �2� 	��Ƴ� 	����)� 	��F�u� 	��        Ƴس 	����"� 	��"�'� P'�)� uF�\� 	��\�p� P        �"� RF�X� R        "�'� P'�)� u\�p� P        �"� P        F�X� R        E�u� u��� u�        E�u� 	���� 	��        E�k� 	��k�u� P��� 	����� P        \�k� R��� R        k�u� P��� P        h�k� P        ��� R        ��� ud��� t`���� ud��� ud��-� ud�-�0� t`�        ߰� 2�        ߰� u$        ߰� u$        ��� ud��� t`��-� ud�-�0� t`�        ��� uc��� t_��-� uc�-�0� t_�        ��� P�"� P        �a� uD        �� ud�� � P �$� ud�$�+� P+�.� t .�1� t1�5� t5�a� ud�        V�a� ud�        ���� u����� P���� u�        *�q� u���� u�[�g� u�        1�C� P��� P        =�C� 1�        ��� P        J�q� u���� u�[�g� u�        J�M� u�M�V� PV�q� u���� u�[�g� u�        ��ö u�ö˶ P˶� u�[�g� u�        ���� uc����� R���� uc�        ���� P        ��,� �         ��,� �        ��� Q�,� �        ��� P�,� �        ��� 2�        ��� �        ���� �        (�+� P+�F� WF�P� UP��� W���� U��� W��� U�� W�6� U6�V� WV��� U���� W��ļ U        (�F� 1�F��� QĹ� Q?�R� QR�X� U���� Q��� Q$�@� Q@�[� �E�� Q�*� �E*�6� Q��ļ Q        (�F� 1�F�|� �D���� �D�� �D�4� S4�G� 0�V��� �D���� 0���ļ �D        ;��� R)�L� R��� R$�@� R@�[� �F��ļ R        B�ӹ S?�|� S���� S�� SV��� S��ļ S        B�R� 0�R�v� P���� 0���� P��� 0���� P�G� 0�V��� 0����� P��ļ 0�        B�F� 0�F�s� V��� V��� V��� V�G� VV�ļ V        �� P��� ��ļ �        ��� P        ]�L� ������ ����� ���G� ��V��� ����ļ ��        ]�L� ������ ����� ���G� ��V��� ����ļ ��        ]�L� 	������ 	����� 	���G� 	��V��� 	����ļ 	��        ]�t� 	��t��� ���� 	����� P�� �$�A� 	��A�[� P[�q� 	����ļ �        ��� P$�@� P        ��� P�� �A�[� P        ���� W        8�@� P        A�[� P        t��� ������ ������ ������ ������ �X�  ��� �W�  �� ���$� �+�  q��� ������ �+�  V�q� ��q��� �X�  ��ļ ��        t��� ��  ���� �N�  ���� �$�  ���� �!�  ���� �N�  ���� �$�  ��� ��  �$� �!�  [�q� ��  q��� �!�  V��� �N�  ���� �$�  ��ļ �!�          t�L� ������ ����$� ��[��� ���G� ��V��� ����ļ ��        t�L� 	������ 	����$� 	��[��� 	���G� 	��V��� 	����ļ 	��        t��� 	������ 	������ P��� 	��[�q� 	��V�q� 	��q��� P        ���� PV�p� P        ���� P���� �q��� P        ���� W        h�p� P        q��� P        ��L� ���$� ��q��� ���G� ������ ����ļ ��        ��L� 	���$� 	��q��� 	���G� 	������ 	����ļ 	��        ���� 	���� 	���$� Pq��� 	������ P��ļ 	��        �$� Wq��� W        �$� P���� P        �� P        ���� W        ���� P        ��L� ���*� ��         �� P�� P        �� 1�        �� P        ��� 2�        ��� �        �	� P	��� uP���� uP��x� uP���� uP��&� uP@�\� uPk�n� uPw��� uP        �	� p� �	��� uP#J����� uP#J���x� uP#J����� uP#J���&� uP#J�@�\� uP#J�k�n� uP#J�w��� uP#J�        �G� 0�G�r� Pr��� SU�\� P���� 	���� P���� P���� S���� P���� S���� S���� P���� S���� P���� S@�K� 0�K�M� PM�R� Sk�w� S        ���� w @)����� w @)����� w @)���#� w @)�@�U� w @)�k��� w @)�        �ʽ uH���� uH��+� uH@�a� uHk��� uH        ,�5� P5��� uO���� 1���� uO��� 0����� 1���� uO�� �G��� uO���� 0����� uO��� 0��Z� uOZ��� 0����� uO��x� 0�x��� 1���+� 0�+�=� uO=�@� �G@�K� PK�R� uOR��� 0�        ,�J� 0�N��� u����� u���+� u�@�K� 0�K�a� u�k��� u�        ���� 0���ʽ uN���� 0���3� uN:��� uN���� 1����� uN��+� uNR�Y� uNk�w� uNw��� 1�        ���� 0���ʽ uD��R� uD��� uD�� ����� uD��� uD��� uD\�k� uD�t� uDx�� uD���� uD	�5� uD�Z� uD���� 0���/� uD:��� uD��=� uD=�@� ��R�w� uD        ʽ� uT�� �L��� uT���� uT+�=� uT=�@� �La�k� uT���� uT        ٽ�� 0���о S�q� Sq��� 0���� 0��� S2�Z� SZ��� 0�a�k� 0�        ٽ� 0��¾ W�q� Wq��� 0����� W��� W�� P�2� W2�D� PD�G� WZ��� Wa�k� W        ٽ�� 	������ 	��+�@� 	��a�k� 	��        �� P�� 
��uH��� 
���@��׿ 
��uH�׿ٿ p uH�ٿf� 
��uH�f�h� r uH�h��� 
��uH����� 
��uH�+�=� 
��uH�=�@� 
���@�a�k� 
��uH�        �� 0��о V�q� Vq��� 0���� V�� R�v� Vv�x� Qx��� V��M� VZ��� Va�k� V        �� 0�q��� 0�M�x� P���� P���� r rr@*( �        �� W�� u@�� uP#N��� �H#N��q� uP#N�q��� W���� u@���� uP#N����� u@��Z� uP#N�Z��� u@+�=� uP#N�=�@� �H#N�a�k� u@        ܼG� SG��� u ���� u @�B� SB�R� u         ��� W��#� s        �� u�� � V �� u��� ���q� u�q��� V���� u����� V���� u���+� V+�=� u�=�@� ��@�a� Va�k� u�k��� V���� u�        �� u��#� P#�5� u�5�=� P=�� u��� ���=� u�=�@� ��@��� u�        2�5� u�5�=� P=��� u����� u���+� u�K�a� u�k��� u�        o��� u����� u�        ���� u����� u�        ���� u����� P���� u����� u�        ʽ� ud��� �\���� ud����� ud�+�=� ud�=�@� �\�a�k� ud����� ud�        ӽٽ ud���� ud        U�\� P���� 	��        ��� uT���� uT��� uT        ��� uP#N����� uP#N���� uP#N�        �w� u���� u\�v� u        �8� 	��8��� S��ÿ 	��ÿ
� S\�k� 	��k��� S        ��Ϳ u\�k� u        ��Ϳ uP#N�\�k� uP#N�        ��Ϳ uT\�k� uT        8��� Sÿ
� Sf��� S        J�R� u���� u�        R�w� Pk�x� P        ^�w� 1�        k�x� P        k�w� u����� u�        k�w� u����� u�        k��� 	������ 	��        k�z� 	��z��� P���� u��� 	������ 	������ P        k�z� P���� P        z��� P���� u���� P        w�z� R        ���� P        ���� �֓  ���� u�
�� u��,� �ϔ  :�R� u�R�\� �%�  ���� u����� �%�  ��� �ϔ          ���� �  ���� �Ŕ  ���� �  ��
� �  
�$� �Ŕ  $�:� �  :�\� ��  ���� ��  ��� �Ŕ          ���� u���� u�        ���� 	����\� 	������ 	����� 	��        ���� 	����� 	���$� P���� 	����� P        �� R���� R        �$� P$�,� u��� P        �� P        ���� R        ��� u��� P�� u�        0�x� �{�  ���� �{�          0�x� uT���� uT        0�x� u@���� u@        �%� P%�&� t &�*� t*�5� uD        �%� ud�%�*� P*�:� ud�        x�� u����� u�        ��� P:�H� P        ���� 1�        :�H� P        ���� u�V�f� u�        ���� u�V�f� u�        ���� 	��V��� 	��        ���� 	������ P���� u���� 	��V�|� 	��|��� P        ���� PZ�x� P        ���� P���� u|��� P        ���� R        f�x� P        ���� �]�  ���� u����� u��	� �V�  l��� �V�          ��� �"�  ���� �%�  ���� �L�  ���� �"�  ���� �%�  ��	� �L�  Z��� �L�          ���� u����� u�        ��� 	������ 	����	� 	��Z��� 	��        ���� 	����� 	���� P�	� uZ�l� 	��l��� P        ��� RZ�h� R        �� P�	� ul��� P        ��� P        Z�h� R        ,�\� u����� u�        ,�\� 	������ 	��        ,�R� 	��R�\� P���� 	������ P        C�R� R���� R        R�\� P���� P        O�R� P        ���� R        ��� ud��� �\��q� ud��Z� ud�+�=� ud�=�@� �\�        ־ܾ 2�        ־ܾ u$        ־ܾ u$        �� ud��� �\�+�=� ud�=�@� �\�        �� uc��� �[�+�=� uc�=�@� �[�        ��� P+�2� P        �a� uD        �� ud�� � P �$� ud�$�+� P+�.� t .�1� t1�5� t5�a� ud�        S�a� ud�        ���� u����� P���� u�        :��� u���� u�k�w� u�        A�S� P��� P        M�S� 1�        ��� P        Z��� u����� u�k�w� u�        Z�]� u�]�f� Pf��� u����� u�k�w� u�        ���� u����� P���� u�k�w� u�        ���� uc����� R���� uc�        ���� P        �<� �         �<� �        �/� Q/�<� �        �/� P/�<� �        ���� P��W� uP!�c� uP&��� uP�J� uPO��� uP���� uP���� uP��� uP        ���� p� ���W� uP#J�!�c� uP#J�&��� uP#J��J� uP#J�O��� uP#J����� uP#J����� uP#J���� uP#J�        ���� 0���� P�A� S���� P|��� 	������ P!�<� P<�E� SE�^� P^�c� S&�<� S<�B� PB�I� S\�i� Pi�x� S���� 0����� P���� S���� S        ��W� w @)�!�c� w @)�&�C� w @)�O��� w @)����� w @)���� w @)�        ��j� uH!�c� uH&��� uH���� uH��	� uH        ���� P��A� uOA�W� 1����� uO��=� 0�=�C� 1�C��� uO���� �G��.� uO7�!� 0�!�c� uOc��� 0����� uO��� 0�&�I� uOI��� 0���� 1���� 0����� uO���� �G���� P���� uO��� 0�        ���� 0���W� uL!�c� uL&��� uL���� 0����� uL��� uL        A�W� 0�W�j� uNI�Z� 0�Z��� uN�� � uN �?� 1�?�G� uNO��� uN���� uN���� uN��� 1�        A�W� 0�W�j� uD���� uD=��� uD���� ����.� uD7�� uD���� uD���� uD���� uD �� uDT�l� uD���� uD���� uDI�Z� 0�Z��� uD��$� uD?��� uD���� ������ uD        j��� uT���� �L��!� uTc�&� uT���� uT���� �L���� uT�.� uT        y�C� 0�C��� S��� S�!� 0�c��� 0����� S��� 0����� 0�        y��� 0���a� W��� W�.� 0�7�!� Wc��� W���� P���� W���� P���� W��� W���� W        y�!� 	��c�� 	������ 	������ 	��        ���� P���� u@���� ����!� u@c�� u@���� u@���� ������ u@        ���� 0���p� V��� V�.� 0�7�{� V���� V �!� Vc��� V��� V���� V        ���� 0��.� 0��� � PT�l� P        ���� W���� u����� uP#N����� �H#N���� uP#N��$� W$�.� u�.��� uP#N���!� u�c��� uP#N���� u����� uP#N����� �H#N����� u�        |��� S��0� u !�c� u ���� S���� u         ���� W���� s        ���� u����� V���� u����� ����� u��"� V"�!� u�!�c� Vc�� u���� V���� u����� ������ V���� u���� V�.� u�        ���� u����� P���� u����� P���� u����� ������ u����� ����.� u�        ���� u����� P��A� u�!�c� u�&��� u����� u���� u�        �A� u�&�I� u�        )�A� u�&�I� u�        )�,� u�,�5� P5�A� u�&�I� u�        j��� ud����� �\���!� ud�c�&� ud����� ud����� �\����� ud��.� ud�        s�y� ud�� ud        ���� P|��� 	��        ��=� uT7��� uTc��� uT        ��=� uP#N�7��� uP#N�c��� uP#N�        ��� u7��� u��� u        ���� 	����)� S7�c� 	��c��� S���� 	����Q� S        7�l� u���� u        7�l� uP#N����� uP#N�        7�l� uT���� uT        ��)� Sc��� S��Q� S        ���� u����� u�        ��� P��� P        ��� 1�        ��� P        
�� u��*� u�        
�� u��*� u�        
�5� 	���Q� 	��        
�� 	���+� P+�5� u���� 	���<� 	��<�Q� P        
�� P�8� P        �+� P+�5� u<�Q� P        �� R        *�8� P        �)� �?�  )�5� u����� u����� �8�  ���� u����� �  Q�l� u�l�|� �  |��� �8�          �)� ��  )�5� �.�  5�=� ��  ���� ��  ���� �.�  ���� ��  ���� �  Q�|� �  c��� �.�          �5� u����� u�        �=� 	������ 	��Q��� 	��c��� 	��        �5� 	������ 	������ Pc�|� 	��|��� P        ���� Rc�x� R        ���� P���� u|��� P        ���� P        c�x� R        ���� u����� P���� u�        �� � ��  T�l� ��          �� � uTT�l� uT        �� � u�T�l� u�        ���� P���� t ���� t���� uD        ���� ud����� P���� ud�         �� u�h�l� u�        �,� R���� R        �,� 1�        ���� R         �,� u����� u�         �,� u����� u�         �G� 	����!� 	��         �/� 	��/�A� PA�G� ul��� 	����� 	���!� P         �/� R��� R        /�A� PA�G� u�!� P        ,�/� P        ��� R        5�?� �Ƨ  ?�G� u����� u����� �  ��� �          ���� �  5�?� �  ?�G� �  G�T� �  l��� �  ���� �  ��� �          5�G� u�l��� u�        ���� 	��5�T� 	��l��� 	����� 	��        5�G� 	��l��� 	������ P���� u���� 	���� � P        ���� R���� R        ���� P���� u�� � P        ���� P        ���� R        ���� u�Q��� u�        ���� 	��Q��� 	��        ���� 	������ PQ�l� 	��l�|� P        ���� RQ�h� R        ���� Pl�|� P        ���� P        Q�h� R        C��� ud����� �\���� ud����� ud����� ud����� �\�        v�|� 2�        v�|� u$        v�|� u$        ���� ud����� �\����� ud����� �\�        ���� uc����� �[����� uc����� �[�        ���� P���� P        ��� uD        ���� ud����� P���� ud����� P���� t ���� t���� t��� ud�        ��� ud�        &�3� u�3�;� P;�I� u�        ��� u�O��� u����� u�        ���� Px��� P        ���� 1�        x��� P        ��� u�O�x� u����� u�        ���� u����� P��� u�O�x� u����� u�        O�S� u�S�[� P[�x� u����� u�        � � uc� �$� R$�.� uc�        �$� P        ���� �         ���� �        ���� Q���� �        ���� P���� �        �)� P)��� uP���� uP��x� uP���� uP��&� uP@�\� uPk�n� uPw��� uP        �)� p� �)��� uP#J����� uP#J���x� uP#J����� uP#J���&� uP#J�@�\� uP#J�k�n� uP#J�w��� uP#J�        �g� 0�g��� P���� Si�p� P��� 	���"� P���� P���� S���� P���� S���� S���� P���� S���� P���� S@�K� 0�K�M� PM�R� Sk�w� S        ��� w @)����� w @)����� w @)���#� w @)�@�U� w @)�k��� w @)�        4��� uH���� uH��+� uH@�a� uHk��� uH        L�U� PU��� uO���� 1��6� uO6��� 0����� 1���"� uO"�%� �G%��� uO���� 0����� uO��� 0��Y� uOY��� 0����� uO��x� 0�x��� 1���+� 0�+�=� uO=�@� tK@�K� PK�R� uOR��� 0�        L�j� 0�n��� uL���� uL��+� uL@�K� 0�K�a� uLk��� uL        ���� 0����� uN���� 0���3� uN:��� uN���� 1����� uN��+� uNR�Y� uNk�w� uNw��� 1�        ���� 0����� uD�q� uD��"� uD"�%� ��%��� uD���� uD�� uDp�{� uD"�|� uD���� uD���� uD�E� uD�Y� uD���� 0���/� uD:��� uD��=� uD=�@� t@R�w� uD        ��"� uT"�%� �L%��� uT���� uT+�=� uT=�@� tPa�k� uT���� uT        ���� 0���� S%��� S���� 0���� 0��Y� SY��� 0�a�k� 0�        ��6� 0�6��� W%��� W���� 0����� W��&� W&�)� P)�@� W@�D� PD�G� WY��� Wa�k� W        ���� 	������ 	��+�@� 	��a�k� 	��        �	� P	�"� u@"�%� ��%��� u@���� u@+�=� u@=�@� t�a�k� u@        �6� 0�6��� V%��� V���� 0����� V�~� V���� V��M� VY��� Va�k� V        �6� 0����� 0�]��� P���� P        �"� W"�6� u�6�"� uP#N�"�%� �H#N�%��� uP#N����� W���� u���� uP#N���� u���Y� uP#N�Y��� u�+�=� uP#N�=�@� tL#N�a�k� u�        ��g� Sg��� u ���� u @�B� SB�R� u         �� W�C� s        4�:� u�:� � V �"� u�"�%� ��%��� u����� V���� u����� V���� u���+� V+�=� u�=�@� t�@�a� Va�k� u�k��� V���� u�        4�7� u�7�C� PC�U� u�U�]� P]�"� u�"�%� ��%�=� u�=�@� t�@��� u�        R�U� u�U�]� P]��� u����� u���+� u�K�a� u�k��� u�        ���� u����� u�        ���� u����� u�        ���� u����� P���� u����� u�        ��"� ud�"�%� �\�%��� ud����� ud�+�=� ud�=�@� t`�a�k� ud����� ud�        ���� ud���� ud        i�p� P��� 	��        6��� uT��� uT��� uT        6��� uP#N���� uP#N���� uP#N�        6��� u��� up��� u        6�X� 	��X��� S���� 	����"� Sp�{� 	��{��� S        ���� up�{� u        ���� uP#N�p�{� uP#N�        ���� uTp�{� uT        X��� S��"� Sv��� S        i�q� u��� u�        q��� P{��� P        }��� 1�        {��� P        ���� u����� u�        ���� u����� u�        ���� 	������ 	��        ���� 	������ P���� u�(� 	������ 	������ P        ���� P���� P        ���� P���� u���� P        ���� R        ���� P        ���� �  ���� u�"�(� u�7�D� �  R�f� u�f�p� ���  ���� u����� ���  ��� �          ���� �p�  ���� �  ���� �m�  �"� �p�  "�<� �  <�R� �m�  R�p� ��  ���� ��  ��� �          ���� u��(� u�        ���� 	���p� 	����� 	����� 	��        ���� 	���7� 	��7�<� P���� 	����� P        (�7� R���� R        7�<� P<�D� u��� P        4�7� P        ���� R        �� u��� P�"� u�        @��� �M�  ���� �M�          @��� uT���� uT        @��� u����� u�        +�5� P5�6� t 6�:� t:�E� uD        +�5� ud�5�:� P:�J� ud�        ���� u����� u�        ���� RJ�X� R        ���� 1�        J�X� R        ���� u�f�v� u�        ���� u�f�v� u�        ���� 	��f��� 	��        ���� 	������ P���� u��� 	��f��� 	������ P        ���� Rj��� R        ���� P���� u���� P        ���� P        v��� R        ���� �/�  ���� u��� u��� �(�  l��� �(�          �"� ���  ���� ���  ���� ��  ���� ���  ��� ���  �� ��  Y��� ��          ���� u���� u�        �"� 	������ 	����� 	��Y��� 	��        ���� 	����� 	���� P�� uY�l� 	��l��� P        �� RY�h� R        �� P�� ul��� P        �� P        Y�h� R        D�p� u���� u�        D�p� 	����� 	��        D�f� 	��f�p� P���� 	������ P        [�f� R���� R        f�p� P���� P        c�f� P        ���� R        ��"� ud�"�%� �\�%��� ud��Y� ud�+�=� ud�=�@� t`�        ���� 2�        ���� u$        ���� u$        �"� ud�"�%� �\�+�=� ud�=�@� t`�        �"� uc�"�%� �[�+�=� uc�=�@� t_�        �� P+�2� P        %��� uD        %�;� ud�;�@� P@�D� ud�D�K� PK�N� t N�Q� tQ�U� tU��� ud�        s��� ud�        ���� u����� P���� u�        :��� u���� u�k�w� u�        A�S� P��� P        M�S� 1�        ��� P        Z��� u����� u�k�w� u�        Z�]� u�]�f� Pf��� u����� u�k�w� u�        ���� u����� P���� u�k�w� u�        ���� uc����� R���� uc�        ���� P        ��H� �L�P� P�R�        �Y� WY�\� �#        �� w 	���� R�Y� w 	��Y�\�
 �#	��        7�W� SW�\� �        7�Y� WY�\� �#        7�B� s        }��� �         }��� �        }��� Q���� �        }��� P���� �        ���� P���� V��6� V^�6� V��0� VB�a� Vv��� V        ���� p� ����� v� ���6� v� �^�6� v� ���0� v� �B�a� v� �v��� v� �        ��X� 0�X�z� Pz��� S���� P4�@� P���� P���� 	������ P���� S���� P��� S�� S�"� P"�� S�+� P+�0� SB�a� Sv��� 0����� P���� S���� P���� S        � � p @)� ��� uH@)���� uH@)��0� uH@)�B�a� uH@)�v��� uH@)����� uH@)�        &��� uP��� uP�0� uPB�a� uPv��� uP���� uP        >�G� PG��� u����� 1�5�R� u�R�}� 0�}��� 1����� u����� ������ 0���}� u���q� 0�q��� u����� 0���� u��6� 0�6��� u����� 0��%� u�%��� 0����� 1���0� 0�0�B� u�B�a� 0�a�s� u�s�v� ��v��� P���� u����� 0�        >�X� 0�\��� u���� u��0� u�B�a� u�v��� 0����� u����� u�        ���� 0����� u�%�0� 0�0��� u����� u����� 1���� u�	�0� u�B�a� u����� u����� u����� 1�        ���� 0����� u�5� � u�&�1� u�}��� u����� ����}� u����� u���� u�q��� u����� u�6�@� u����� u�6��� u�%�0� 0�0�� u����� u���s� u�s�v� ������ u�        ��� uH��� uH        ���� 0����� S���� 0���^� S^��� 0��6� 0�6��� S���� 0�0�B� S���� 0�        ��R� 0�R��� W��^� W^�}� 0���q� Wq��� 0����� W�F� WF�M� PM�q� Wq��� P���� W0�B� W���� W         �� u�        #�R� u��R�R���
 u��u������
 ��������^�
 u��u��^�}� u��R�}�q�
 u��u��q��� u��R�����
 u��u�����
 u��u��0�B�
 u��u��a�s�
 u��u��s�v�
 ����������
 u��u��        #�R�
 �        R��� uP��#� uP&�1� uP}��� uP���� �H��^� uP^�}�
 �        ���� uP��� uPq���
 �        ���� uP���� uP6�@� uP���� uP���� uP6��� uP0�B� uPa�s� uPs�v� �H���� uP        #�R� 0����� P���� R���� u�^�}� 0����� Rq��� 0�        &�*� P*�}� u�}��� v� ����� u���6� v� �^�}� u�}��� v� ����� u����� v� ��6� v� ����� u����� u�        ��X� SX��� u ��� u v�x� Sx��� u         ��0� s        &�,� u�,��� W���� u����� ������ u���� W�� u��0� W0�B� u�B�a� Wa�s� u�s�v� ��v��� W���� u����� W���� u�        &�)� u�)�5� P5�G� u�G�O� PO��� u����� ����s� u�s�v� ��v��� u�        D�G� u�G�O� PO��� u���� u��0� u�B�a� u����� u����� u�        w��� u��%� u�        ���� u��%� u�        ���� u����� P���� u��%� u�        ���� ud����� �\����� ud��� ud�0�B� ud�a�s� ud�s�v� �\����� ud����� ud�        ���� ud���� ud        x�&� ��  ���� ��  ���� ��          x�&� uH���� uH���� uH        x�&� u����� u����� u�        ��� P�� t �
� t
�� u�        ��� ud��
� P
�� ud�        &�1� u����� u�        1�V� P�(� P        =�V� 1�        �(� P        J�V� u�6�J� u�        J�V� u�6�J� u�        J�u� 	��6�q� 	��        J�Y� 	��Y�k� Pk�u� u���� 	��6�\� 	��\�q� P        J�Y� P>�X� P        Y�k� Pk�u� u\�q� P        V�Y� R        J�X� P        _�i� �c�  i�u� u����� u����� �\�  ���� �\�          _�i� �+�  i�u� �R�  u�}� �(�  ���� �+�  ���� �R�  ���� �(�  ���� �R�          _�u� u����� u�        _�}� 	������ 	������ 	��        _�u� 	������ 	������ P���� 	������ P        ���� R���� R        ���� P���� u���� P        ���� P        ���� R        ���� u����� P���� u�        4�@� P���� P���� 	��        ���� uH6�@� uH        ���� v� ��6� v� �        ���� u6�@� u        ���� 	������ u�6�o� 	������ u�)�>� 	��        @�o� u)�>� u        @�o� v� �)�>� v� �        @�o� uH)�>� uH        ���� Pj�o� P���� P9�>� P        ���� u����� u�        ���� P>�H� P        ���� 1�        >�H� P        ���� u�V�f� u�        ���� u�V�f� u�        ��� 	��V��� 	��        ��� 	���� P�� u��� 	��V�|� 	��|��� P        ��� PZ�x� P        �� P�� u|��� P        ��� R        f�x� P        �� ���  �� u�/�6� u�o�� u���� ��  
�� u��)� ���  ���� u����� ��  �6� ���          �� ��  �� ���  �/� ��  /�@� ��  o��� ��  ��
� ��  
�)� ���  ���� ��  �6� ���          �� u���� u�        �@� 	��o��� 	����)� 	������ 	���6� 	��        �� 	����� 	���$� P$�)� u�� 	���1� P        �� R�� R        �$� P$�)� u�1� P        �� P        �� R        !�@� u�o��� u����� u�        !�@� 	��o��� 	������ 	��        !�6� 	��o�� 	����� P���� 	������ P        o�� R���� R        ��� P���� P        |�� P        ���� R        ���� ud����� �\���^� ud�6��� ud�0�B� ud�a�s� ud�s�v� �\�        ���� 2�        ���� u$        ���� u$        ���� ud����� �\�a�s� ud�s�v� �\�        ���� uc����� �[�a�s� uc�s�v� �[�        ���� Pa�h� P        ��N� u�        ��� ud��� P�� ud��"� P"�N� ud�        @�N� ud�        �� u��� P�%� u�        ���� u�	�0� u�B�a� u����� u�        ���� PB�X� P        ���� 1�        B�X� P        ���� u�	�0� u����� u�        ���� u����� P���� u�	�0� u����� u�        	�� u��� P�0� u����� u�        ���� uc����� R���� uc�        ���� P        =�l� �         =�l� �        =�_� Q_�l� �        =�_� P_�l� �        ���� P���� u@A��� u@U��� u@��� u@�,� u@        ���� p� ����� u@#J�A��� u@#J�U��� u@#J���� u@#J��,� u@#J�        ��� 0��?� P?�n� S���� P,�6� 	������ PA�\� P\�e� Se�~� P~��� Sv��� S���� P���� S���� P���� S���� 0����� P���� S�� P�� S        ���� p @)����� uP@)�A��� uP@)�v��� uP@)����� uP@)�        ���� VA��� VU��� V��� V�'� V        ��� P�n� u�n��� 1����� u����� 0����� 1��� � u� �� t���� u���A� 0�A��� u����� 0���+� u�+�U� 0�v��� u���@� 0�@�P� 1�P��� 0����� u����� t����� P���� u���,� 0�        ��� 0���� u�A��� u�v��� u����� 0���� u��,� u�        n��� 0����� u����� 0���� u��[� u�[�y� 1�y��� u����� u����� u��� u��,� 1�        n��� 0����� u���H� u��� � u� �� t���� u���.� u�4�<� u����� u�6�M� u�S�^� u���� u����� u���+� u����� 0���� u��_� u�y��� u����� t���� u�        ���� uDU�v� uD        ���� 0����� S�n� Sn�A� 0����� 0����� S+�U� 0��� 0�        ���� 0���H� uH���� uH�n� uHn��� 0���<� uH���� uH6�^� uH��� uH���� uH��� uH�� uH        ��A�
 �����������U�
 �������������
 �����������
 ���������        ���� u��R��� �
 u��u�� ��
 t��t���n�
 u��u��n��� u��R���A�
 u��u����U�
 u��u������
 u��u������
 t��t����
 u��u��        ����
 �        ��H� uP�� � uP �� tL�n� uPn���
 �        ���� uP��(� P�R�4�<� uP���� P�R�6�S� P�R�S�^� uP��9� uP?�b� P�R�b�� uP���� uP��+� uP���� uP���� tL�� uP        ���� 0�n��� 0�6�G� VG�P� uP ����� P��6� Q6�b� Vb�� Q        ���� V�� � u@#N� �� t�#N��n� u@#N�n��� V��6� u@#N�6�A� u���+� u@#N�+�U� u����� u@#N����� t�#N��� u�        ��� S�]� u A��� u ���� S���� u         ���� s        ���� u����� W�� � u� �� t��n� u�n��� W��A� u�A��� W��U� u�U��� W���� u����� t���� W�� u��,� W,�L� u�        ���� u����� P��� u��
� P
� � u� �� t���� u����� t���L� u�        ��� u��
� P
�n� u�A��� u�v��� u���� u��,� u�        <�n� u�v��� u�        V�n� u�v��� u�        V�Y� u�Y�b� Pb�n� u�v��� u�        �� � ud� �� t`��A� ud���v� ud����� ud����� t`��� ud�,�L� ud�        ���� udU�i� ud        ���� P,�6� 	��        ���� uD��6� uD���� uD        ���� u@#N���6� u@#N����� u@#N�        ��m� u��<� u���� u        ��� 	���H� Q���� 	������ Q��%� V%�1� uP ����� V        ���� u        ���� u@#N�        ���� uD        ���� Q        @�H� u�4�<� u�        H�m� P���� P        T�m� 1�        ���� P        a�m� u����� u�        a�m� u����� u�        a��� 	����� 	��        a�p� 	��p��� P���� u<�X� 	������ 	����� P        a�p� P���� P        p��� P���� u��� P        m�p� R        ���� P        v��� ���  ���� u�R�X� u�g�t� ���  ���� u����� �$�  �� u��,� �$�  ���� ���          v��� ��  ���� ���  ���� ��  <�R� ��  R�l� ���  l��� ��  ���� ��  �,� ��  ���� ���          v��� u�<�X� u�        v��� 	��<��� 	���6� 	������ 	��        v��� 	��<�g� 	��g�l� P���� 	������ P        X�g� R���� R        g�l� Pl�t� u���� P        d�g� P        ���� R        6�S� �z�  ��� �z�          6�S� uD��� uD        6�S� u���� u�        ���� P���� t ���� t���� u�        ���� ud����� P���� ud�        S�^� u�w�� u�        ^��� P���� P        j��� 1�        ���� P        w��� u��� u�        w��� u��� u�        w��� 	���A� 	��        w��� 	������ P���� u��� 	���,� 	��,�A� P        w��� P�(� P        ���� P���� u,�A� P        ���� R        �(� P        ���� ��  ���� u����� u����� ��  <�U� ��          ���� ���  ���� ��  ���� ���  ��� ���  ���� ��  +�U� ��          ���� u���� u�        ���� 	����� 	��+�U� 	��        ���� 	����� 	������ P���� u+�<� 	��<�P� P        ���� R+�8� R        ���� P���� u<�P� P        ���� P        +�8� R        ���� u����� P���� u�        t��� u��6� u�        t��� 	���6� 	��        t��� 	������ P�� 	���,� P        ���� R�� R        ���� P�,� P        ���� P        �� R        �� � ud� �� t`��n� ud���+� ud����� ud����� t`�        ���� 2�        ���� u$        ���� u$        �� � ud� �� t`����� ud����� t`�        �� � uc� �� t_����� uc����� t_�        ���� P���� P        �^� u�        �� ud��F� VF�^� ud�        P�^� ud�        v��� u����� P���� u�        �P� u����� u��� u�        �%� P���� P        �%� 1�        ���� P        ,�P� u����� u��� u�        ,�/� u�/�8� P8�P� u����� u��� u�        ���� u����� P���� u��� u�        4�>� uc�>�B� RB�L� uc�        4�B� P        ���� �         ���� �        ���� Q���� �        ���� P���� �         �w� � ��� �          �7� 0�7�P� P        d��� R        d��� 0�        d��� �`�        d��� S        d��� U        ���� ��}�        ���� 1�        ���� ��}�        ���� S        ���� U         �j� � ���� �          �7� 0�7�P� P        ]��� R        ]��� �`�        ]��� S        ]��� U        ��@� S        [��� S        ��@� S        9�=� t J��� t %�)� t 6��� t ���� t ���� t A�E� t b�f� t ���� t         A�E� t         ���� t ��� t ���� t         ���� t         %�)� t 6��� t ���� t ���� t b�f� t ���� t         ���� t         ���� t ���� t b�f� t         b�f� t         �-� 
  �        !�-� 1�        ���� P        ��� �         ��� P        ^�m� Sm�o� Po��� S        i�h� uw�o��� uw�        i�h� 1�o��� 1�        o��� Ro�w� R        ���� S���� u���� sd����� uL����� tL����� S�� � u �� sd�        ���� u���� sd����� uL����� tL�        ���� S�� � u �� sd�        0�C� � L�[� R_�r� R���� R        0�C� �L�[� Q_�y� Q���� Q        ?�C� PC�s� � #���� � #        ���� R        L�[� R���� R        S�[� P���� P        U�[� S���� S        i�r� R        ���� S��� u�� t�R� SR�U� uU�V� tV�i� S        0�V� 	��        0�R� SR�U� uU�V� t        0�R� s,80.�R�U� u#,80.�U�V� t#,80.�        N�V� 0�        N�R� SR�U� uU�V� t        0�V� P        ���� S���� u���� t��� S�� u�� t        ��� 	��        ��� S�� u�� t        ��� s,80.��� u#,80.��� t#,80.�        ��� 0�        ��� S�� u�� t        ��� P         �%� �         0�5� �         G�g� 0�g��� W���� P��� W�� P�=� W=�\� 0�        g��� P���� P���� P���� PK�\� P        V��� S���� � ��� S�� � �\� S        b�e� P        x��� V��� V�=� V        ���� P        }��� V        }��� Q        }��� U        ���� S        ���� S�=� S        ���� 	���=� 	��        ���� S        ���� S        ���� P        ���� P        )�8� P        ���� 1�        �=� S        ���� P���� P        ��� U�=� U        ��� P        ���� 1�        ���� P        ��� U        ��� ��          `��� � ���� R        `��� 	������ P���� 	������ P        j��� �         j��� � # 80.�        x�}� Q        x�}� � #        x�}� � #        x�}� �         ���� � ���� P���� �         ���� P        ���� � # 80.����� p 80.�        ���� � ���� P        ���� � # 80.����� p 80.�        ���� R        ���� p        ���� p        ���� P        ���� P���� � #        ��'� � '�G� Q        ��+� �+�5� P5�<� �<�E� PE�G� �        ��'� 	��'�+� P+�8� 	��8�<� P<�G� 	��        � � � # @0.�        �'� r�        �'� ��          �'� �         �'� 	��        +�<� Q        +�<� 	��        8�<� ��          ��ɀ PɀҀ �P�        ��ɀ RɀҀ �R�        ��ɀ p�ɀҀ �P#�        ���� Q��р s�        b�y� s$�y��� � #$����� s$�        e��� �o����� P���� �o�        e�m� R���� R        ���� �o����� P���� �o�        ���� R        ���� r�        ���� Q���� v�        m�y� Sy��� �         ���� S���� � ��� S        ���� s$����� � #$���� s$�        ��� �o��
� P
�� �o�        ���� R��
� R        ��� �o��
� P
�� �o�        ��
� R        ��
� r�        ��
� Q
�� v�        ���� S���� �         )�K� s�K�e� � #�e��� s�        0�K� s(�K�e� � #(�e��� s(�        3��� �o����� P���� �o�        3�;� Re��� R        e��� �o����� P���� �o�        e��� R        e��� r�        s��� Q���� v�        ;�K� s�K�e� � #�        ���� s���� � #��0� s�        ���� s,���� � #,��0� s,�        ��$� �o�$�*� P*�0� �o�        ���� R�*� R        �$� �o�$�*� P*�0� �o�        �*� R        �*� r�        �*� Q*�0� v�        ���� s���� � #�        Y��� S���� � ���� S        i��� s����� � #����� s�        p��� s(����� � #(����� s(�        s��� �o����� P���� �o�        s�{� R���� R        ���� �o����� P���� �o�        ���� R        ���� r�        ���� Q���� v�        {��� s����� � #�        ���� s,����� P���� s,����� � #,�        ��L� SL�N� � N�p� S        	�L� s�L�N� � #�N�p� s�        �L� s,�L�N� � #,�N�p� s,�        �d� �o�d�j� Pj�p� �o�        �� RN�j� R        N�d� �o�d�j� Pj�p� �o�        N�j� R        N�j� r�        S�j� Qj�p� v�        �L� s�L�N� � #�        .�1� s0�1�?� P?�L� s0�L�N� � #0�        ���� s����� � #���  s�        ���� s0����� � #0���  s0�        ��  �o� 
  P
   �o�        ���� R��
  R        ��  �o� 
  P
   �o�        ��
  R        ��
  r�        ��
  Q
   v�        ���� s����� � #�        I �  S� �  � � �  S        ` �  s�� �  � #�� �  s�        g �  s0�� �  � #0�� �  s0�        j �  �o�� �  P� �  �o�        j r  R� �  R        � �  �o�� �  P� �  �o�        � �  R        � �  r�        � �  Q� �  v�        r �  s�� �  � #�        � �  s4�� �  P� �  s4�� �  � #4�        Y SYZ �         UY s$�YZ � #$�        UY s$YZ � #$        c� u�� u�I u        t� s �� s � s         �� ur��� P�� ur�        �� Q        �� r        �� ut��� P�� ut�        �� P�� ut�        �� u        �� ut��� ut�        �� us��� us�        �� R�� R        �� us��� P�� us�        �� R        �� 	��        �� r�        �� Q�� v�        �� ur��� Q�� ur� ur�        �� P        �� r        �� ut��� P�� ut� ut�        �� P�� ut� ut�        �� u u        � r$� R u#$�        � u        1 ut�        ", us�,0 R01 us�        "0 P        1I u        6@ ut�@D RDN ut�        6D P        Pr � r� P        Zf q 80.�fr � # 80.�r� q 80.�        hn R        hn �         �� � �� S�� �         �� ��� P�R��� P�R�        �� � �� S�� �         �� �         �� ����        �� S�� �         �� P         / �/9 0�9� �         P w 0.�Xi w 0.�in s 80.��� w 0.��� s 80.�        #P q 0.�Xv q 0.��� q 0.�        %W UX� U        %' p r "�'/ R/9 U9P RXv R�� R        #T s$�TX � #$�X� s$��� � #$�        P s Xn s �� s         %T s$�TX � #$�X� s$��� � #$�         P s Xn s �� s         =P U�� U        =I p �"�IP V�� V�� s�� p �"��� ��"�        =P P�� P�� �        =P S�� S�� �         w� U        w� S        �� 0��� Q�� 0��� Q�� 0�        �� p$��� � #$�         � #$� P* � #$�        <| s @0.��� s @0.�x� s @0.��� u# @0.��� t# @0.��� s @0.�        il Pl| s$8�� s$8�� uTx� s$8        i� ���?��� ���?��� ���?�        i| R�� Rx� R        R� s$��� s$��� s$�        x� P�� uT1$�        �� ud��X WXx ud��� W        �� w         �x V�� Q�� V        �x ud��� ud�        �� Q�x uT�� uT         �  �� �           p r "�        x ud��� ud�        x uT�� uT         pt��� pt�        �� uT        �� pt�        �� p uT"�        Cx ud�        Ff uc�fo Pox uc�        Fo R        Rf uc�fo Pox uc�        Ro R        Rx 	��        Ro r�        Uo Qox w�        �� �0  �� �0          �� �  �� �          �� uc��� R�� uc�        �� P        |� S        |� 1�         P; �        - s         : S:; �         , 0�,5 R        ), s$�        L� S�� u�� t� S        �� P�� u�� t�	 u        �� V�� u�� t�� u�� u        �� S�� u�� t�� S�� S        �� 0��� R�� 0�        �� s$�        �� s$�        �� ug��� R�� ug�        �� P        `� Q�� s q ��� R� �Lj ��@H$0)p �80.�y� R�� �L�� �L�� ��@H$0)p �80.��e	 �L        lv Sv� W�� R�e	 �K        z� U�e	 U        �j R�� R�e	 R        Wc Vcj p y� p �e	 p         `c Vcj p y� p �e	 p         �U t Ur �@ry t �� t �	 t �%�X�%"�:	M	 t Q	e	 t         �� t �y �P�� �P�)	 t -	:	 �P:	M	 t Q	e	 t         �j Pjy ��e	 P        �� �P0.��j p 80.��� �P0.��� p 80.��"	 �P0.�"	e	 p 80.�        �� Q        �� P        4 p        * pt "�*/ Q/4 p        4 p        4 P        �	�	 V�W���	G
 V�W��L
�
 V�W��        �	�	 �_        �	�	 �X        �	�	 Q�	-
 QL
c
 Q        �	�	 Q�	-
 r L
�
 r         �	-
 P-
L
 � L
�
 P�
�
 �         �	�	 Q�	-
 r L
�
 r         
L
 1�X
�
 1�        �	-
 R-
L
 �L
�
 R�
�
 �        �	
 u 0.�
-
 r 80.�L
X
 u 0.�X
�
 r 80.�        L
X
 S        L
X
 R        X
o
 r        X
e
 rv "�e
o
 Q        X
o
 r        X
o
 R        �
< v�<> u#�>? t#�?b v�        �
; S;> u>? t?b S        �
> u8!�>? t8!�?b u8!�        �
= W=> u#�>? t#�?b W        $= w$�=> u#,�>? t#,�?b w$�        $' s,        �
> u>? t?b u        | s0�W VWY u#0�YZ t#0�Z� V        �V SVY uYZ tZ� S        �Y u8!�YZ t8!�^p u8!�        � s�X WXY u#�YZ t#�^m Wmp s�        FX w$�XY u#,�YZ t#,�^m w$�mp s,�        FI s,        �Z 8�^p 8�        �Y uYZ t^p u        �y v�y{ u#�{| t#�|� v�        �x Sx{ u{| t|� S        �� u8!�� P{ uT{| tP|� uT�� u8!��� uT�� u8!�        �{ u{| t|� u�� u        �z Wz{ u#�{| t#�|~ W~� s��� W�� s��� W        02 P2{ u{| t|� u�� u        C{ uT{| tP�� uT�� u8!��� uT�� u8!�        Cz Wz{ u#�{| t#��� W�� s��� W        OW 0�W` R        TW w$�        �� s,�        �� ug��� R�� ug�        �� P        �� s�        �{ u{| t|� u        �� v�        �� S        �� s0�� V u#0� t#0�k V        5 S u tk S        f 8�: 8�Rk 8�        f� P� u t: uRk u        p� p 8!��� P� uT tP uT u8!�: uTRc u8!�ck uT        p u t2 uRk u        p W u#� t#� W: s�R^ W^c s�ce Weg s�gi Wik s�        � u t2 uRk u        � uT tP uT u8!�% uTRc u8!�cg uT        � W u#� t#� W% s�R^ W^c s�ce Weg s�        �� 0��� R        �� w$�        % s,�          ug� $ R$% ug�        $ P        %: s�        :R s0�        �� s��� � #��� s�        �� s,��� � #,��� s,�        �� �o��� P�� �o�        �� R�� R        �� �o��� P�� �o�        �� R        �� r�        �� Q�� w�        �� s��� � #�        �� v��� �#�        �� S�� �         4 r�4U u#�`n r�n� u#��� r��� u#�        U u`� u�� u        , s `f s �� s         &) ur�)4 P4D ur�        &4 Q        &+ r        &< ut�<C PCD ut�        =C PCD ut�        =D u        JU ut��� ut�        MU us��� us�        MU R�� R        �� us��� P�� us�        �� R        �� 	��        �� r�        �� Q�� v�        `c ur�cn Qn� ur��� ur�        `n P        `e r        `v ut�v} P}� ut��� ut�        w} P}� ut��� ut�        w� u�� u        �� r,��� R�� u#,�        �� u        �� ut�        �� us��� R�� us�        �� P        �� u        �� ut��� R�� ut�        �� P        / V/0 � #�        ! s(        / V/0 � #�          0� ) R          v$�        ?� v��� u#��� t#��� v�        ?� S�� u�� t�� S        f� u@!��� t@!��� u@!�        f� W�� u#��� t#��� W        �� w$��� u#(��� t#(��� w$�        �� s(        f� u�� t�� u         s,�� V�� u#,��� t#,�� V        U� S�� u�� t� S        |� u@!��� t@!��� u@!�        |� s��� W�� u#��� t#��� W�� s�        �� w$��� u#(��� t#(��� w$��� s(�        �� s(        |� @��� @�        |� u�� t�� u        /� v��  u#�  t#�` v�        /� S�  u  t` S        \~ u@!�~� P�  uT  tP uT
 u@!�
8 uT8` u@!�        \  u  t. uO` u        \� W�  u#�  t#� W s� WO s�O` W        �� P�  u  t. uO` u        �  uT  tP uT
 u@!�
! uTO` u@!�        �� W�  u#�  t#� W! s�O` W        �� 0��� R        �� w$�        ! s(�         ug�  R ! ug�          P        !8 s�        \  u  t` u        8O v�        8O S        lo s,�o} V} u#,�� t#,��� V        �| S| u� t�� S        �� @��� @��� @�        �� P� u� t�� u�� u        �� p @!��# P# uT� tP�� uT�� u@!��� uT�� u@!��� uT        � u� t�� u�� u        �~ W~ u#�� t#��� W�� s��� W�� s��� W�� s��� W�� s�        ; u� t�� u�� u        N uT� tP�� uT�� u@!��� uT�� u@!��� uT        N~ W~ u#�� t#��� W�� s��� W�� s��� W�� s�        Zb 0�bk R        _b w$�        �� s(�        �� ug��� R�� ug�        �� P        �� s�        �� s,�        E s�EH � #�Hp s�        E s(�EH � #(�Hp s(�        d �o�dj Pjp �o�          RHj R        Hd �o�dj Pjp �o�        Hj R        Hj r�        Sj Qjp w�         E s�EH � #�        3F v�FH �#�        3E SEH �         �� r��� u#��� r�� u#�& r�&i u#�        �� u� ui u        �� s �� s ' s         �� ur��� P�� ur�        �� Q        �� r        �� ut��� P�� ut�        �� P�� ut�        �� u        �� ut�  ut�        �� us�  us�        �� R  R          us� P us�          R          	��          r�         Q v�        �� ur��� Q�  ur�:< ur�        �� P        �� r        �� ut��� P�  ut�:< ut�        �� P�  ut�:< ut�        �  u:< u        & r(�&, R,2 u#(�        2 u        <Q ut�        BL us�LP RPQ us�        BP P        Qi u        V` ut�`d Rdn ut�        Vd P        �� V�� � #�        �� s$        �� V�� � #�        �� 0��� R        �� v$�        �� v��� u#��� t#��� v��� u#�        �� S�� u�� t�� S        �� v��� u#��� t#��� v��� u#�        �� v��� u#��� t#��� v��� u#�        �� s��� u#��� t#��� s�        �� v�        �� S        C� u�� t�� u�� u        C� W�� u#��� t#��� W�� W        w� w$��� u#0��� t#0��� w$��� w$�        wz s0        �� s4��� V�� u#4��� t#4�� V        %� D	��� t �� t� D	�        %� S�� u�� t� S        E� P	��� P	�        E� s��� u#��� t#��� s�        r� u�� t�� u        r| s�|� W�� u#��� t#��� W�� s�        �� w$��� u#0��� t#0��� w$��� s0�        �� s0        /2 v�24 u#�45 t#�5z v�z� V�� v�        /1 S14 u45 t5� S        /2 v�24 u#�45 t#�5z v�z� v��� v�        Q2 v�24 u#�45 t#�5z v�z� v��� v�        Q1 s�14 u#�45 t#�5� s�        �� v�        �� S        �4 u45 t5K uM{ u�� u        �4 u45 t5K uMo u�� u        �3 W34 u#�45 t#�5I WIK s�M� s��� W�� s��� W�� s�        �4 u45 t5K uMo u�� u         P4 u45 t5C PCG uMb u�� u        3 W34 u#�45 t#�5G WMb s��� W�� s��� W�� s�         0� R5G 0�        
 w$�        Mb s0�        S] ug�]a Rab ug�        Sa P        bw s�        �� s4��� V�� u#4��� t#4��x V        = D	�=> t >B tBx D	�        � S�� u�� t�x S        5 P	�F P	�^x P	�        5� s��� u#��� t#�� s�F s�^x s�        l� u�� t� u7 u^x u        l� u�� t� u. u^x u        l� W�� u#��� t#�� W s�F s�^e Weg s�gs Wsx s�        �� u�� t� u. u^x u        �� P�� u�� t� u! u^x u        �� W�� u#��� t#�� W! s�^e Weg s�gs Wsx s�        �� 0��� R� 0�        �� w$�        ! s0�         ug�  R ! ug�          P        !6 s�        F^ s4�        �� s�� � #�0 s�        �� s0�� � #0�0 s0�        �$ �o�$* P*0 �o�        �� R* R        $ �o�$* P*0 �o�        * R        * r�        * Q*0 w�        �� s�� � #�        �  v�  �#�        �� S� �         �  v�  �#�        �� s�� � #�        �  v�  �#�        �� S� �         Nt r�t� u#��� r��� u#��� r��) u#�        N� u�� u�) u        Tl s �� s �� s         fi ur�it Pt� ur�        ft Q        fk r        f| ut�|� P�� ut�        }� P�� ut�        }� u        �� ut��� ut�        �� us��� us�        �� R�� R        �� us��� P�� us�        �� R        �� 	��        �� r�        �� Q�� v�        �� ur��� Q�� ur��� ur�        �� P        �� r        �� ut��� P�� ut��� ut�        �� P�� ut��� ut�        �� u�� u        �� r0��� R�� u#0�        �� u        � ut�         us� R us�         P        ) u          ut� $ R$. ut�        $ P        Bo Vop � #�        Oa s,        Oo Vop � #�        O` 0�`i R        ]` v$�        p� � �� r��        �� � #��� r��        �� P�� px�        �� P�  �E   p|�         )  s) /  R/ A  p         P �  8�� �  V� ! u`!'! 8�'!6! u`>!y! 8�y!�! u`�!�! 8��!�! V        f �  W� ! u\!<! W>!d! Wd!e! u#$�e!f! t#$�f!y! W�!�! W        � �  p 3$r "�� �  p3$r "�        � �  0�� ! R        �!�! s��!�! u#�        �!�! s        >!y! 1��!�! 1�        >!b! s�b!e! u#�e!f! t#�f!y! s��!�! s�        >!L! s        "8" S<"f" S        |"�" P�"�" S        �"�" P�"�" S        �"�" 	��        �"�" p��"�" s�        �"�" R�"�" 0��"�" P�"�" r�        �"�" S        P#`# �`#c# �#�c#w# Rw#�# r��#�# r��#�# Q�#�# R�#�# Q�#�# R        �#�# P�#�# P        �#�# 
 @�        �#$ � $a$ Wa$b$ � b$i$ W        �#b$ �b$g$ Pg$i$ �        �#$ R$_$ st1�_$b$
 �<1�b$i$ R        �#F$ RF$I$ r�I$R$ Rb$i$ R        �#$ 1�$$ P$$ 1�$@$ P@$F$ 1�F$b$ Pb$i$ 1�        �#$ 0�$!$ Q!$$$ q�$$($ Qb$i$ 0�        �$�$ u        �$�$ 1��$�$ p 0)��$% 1�%#% p 0)�        �$�$ S�$% s�%+% S        +%I% S        C%U& =��&�& =��&' =�        I%�% S�&' S        g%x% � �  �%�% �!�  &'& �-�  �&�& �-�  �&�& �!�  �&�& � �          g%m% p r "�        m%�% S�&' S        m%{% pt��&' pt�        �&' S        �&' pt�        �&' p s "�        �%�% S        �%U& ;��&�& ;�        �%�% W�&�& W        �%�% �!�  &'& �-�  �&�& �-�  �&�& �!�          �%�% p r "�        �%�% W�&�& W        �%�% pt��&�& pt�        �&�& W        �&�& pt�        �&�& p w "�        �%�% W        �%U& =��&�& =�        �%5& W�&�& W        &'& �-�  �&�& �-�          & & p r "�         &5& W�&�& W         &*& pt��&�& pt�        �&�& W        �&�& pt�        �&�& p w "�        5&U& W        p&�& uP�&�& �H        �&�& *�        �&�& u        �&�& 1�        �$�$ u�&�& u        �$�$ v �&�& v         
'' Q'3' Q        '-' ug�-'3' P3'9' ug�        '3' Q        '3' q�        (( P        �'�' ud��'�' t`�(�( ud�        �'�' V�'�' u`��'�' t\�(�( V        �'�' ud��'�' t`�(�( ud�        (( R        (%( S        (%( W        �'�' u`��'�' t\�%(�( u`�        �'�' u_��'�' t[�%(�( u_�        �'�' Q�'�' uT%(C( uTV(c( Qc(�( uT        V(t( u_�t(�( Q�(�( u_�        V(�( uT        V(�( 	��        V(�( uT#�        c(t( Qt(�( r�        �'�' ud��'�' t`�%(V( ud�        �'�' u`��'�' t\�%(V( u`�        �'�' R�'�' st�%(I( RI(V( st�        %(V( u`�        %(I( RI(V( st�        %(V( 	��        %(I( r�I(V( s|�        3(I( QI(V( w�        �(�( ud��(�( ud�        �(�( u_��(�( u_�        �(�( R�(�( R        �(�( u_��(�( P�(�( u_�        �(�( R        �(�( r�        �(�( Q�(�( w�        �() 0�)) P)') 0�')+) P+)7) 8�7)G) 2�G)W) @�W)}) 0�        �)�) 0��)8* S+*+ S8+:+ S        *%* P        *4* 	��+*+ 	��8+:+ 	��        *%* p�        ** R*4* w�+*+ w�8+:+ w�        K*V* 0�V*�* S�*+ S        o*�* P        o*�* 	���*+ 	��        o*�* p�        r** R*�* w��*+ w�        Z+j+ Sj+k+ � k+�+ S�+�+ �         \+x+ P        k+�+ S�+�+ �         �+�+ R        �+�+ V�+�+ V        �+�+ Q�+�+ w�        �+�+ V        C,I, 0�I,�, R        c,g, Q        c,g, 1�        c,g, q�        �,�, 0��,�, R        �,�, Q        �,�, 1�        �,�, q�        �,�, 0�        -(- P(-P- ud        /'/ V�/�/ V        �-�- R�-�. u�/�/ u�/0 u        �-�- 1�        �-�- �E�        �-�- �E�-�- p�        �-�- P�-. V.A. udA.�. u`#��/�/ u`#��/0 u`#�        �-�- V�-�- s�-�. u\�/�/ u\�/0 u\        .. P.�. V�/�/ V�/0 V        O.Q. PQ.e. se.�. uX�/�/ uX�/0 uX        .. 0�         .L. R        l.�. 0�        �.�. Q        �./ u�/�/ u        �.w/ 1��/�/ 1��/�/ 1�00 1�        �./ u#��/�/ u#�        // P�/�/ P        // 	���/�/ 	��        // p��/�/ p�        // R�/�/ R�/�/ q�        /)/ 0�)/w/ V�/�/ V�/�/ V        O/i/ P        S/i/ P        )/6/ 	��S/w/ 	���/�/ 	���/�/ 	��        S/i/ p�        V/i/ Qi/m/ w��/�/ w��/�/ w�         0a0 � s0�0 �          0i0 �s0�0 �         0e0 �s0�0 �        )0r0 Qs00 Q0�0 �        70F0 1�        70F0 �E�        70D0 �ED0F0 p�        �0�0 ��0�0 S�0�0 s|��0�0 S        �0
1 � 
161 W        �0
1 �
161 S        �0
1 �
161 V        �01 S        �01 1�        �01 s�        J1Y1 1�        J1Y1 �E�        J1W1 �EW1Y1 p�        2!2 � !2%2 pd�        82O2 SO2S2 �         `2u2 �u2�2 U�2�2 U�2�2 u v "��2�2 U        `2y2 0�y2�2 S�2�2 P�2�2 S�2�2 S        �2�2 wp ��2�2 R�2�2 R        y2�2 W�2�2 W        �2�2 �s ��2�2 Q        �2�2 V        �2�2 U        �2�2 P        �2�2 W         33 	��33 P343 	��43?3 P        .3>3 S>3?3 �         1373 R73:3 s:3?3 r�        43>3 S>3?3 �         @3U3 �U3�3 U�3�3 U�3�3 u w "��3�3 U�3�3 R�34 U        @3Y3 0�Y3�3 V�3�3 P�3�3 V�3�3 V�3�3 v��34 V        c3h3 sp �h3j3 R�3�3 R        Y3�3 S�34 S        �3�3 �v ��3�3 Q        �3�3 W        �3�3 P        �3�3 U        �3�3 S        �3�3 P
44 P        w3�3 S�34 S        w3�3 	���34 	��44 P        44 R4
4 s
44 r�        �3�3 �W          4M4 SM4O4 wd�S4p4 Sp4�4 u        55 �        55 �        55 �        55 V55 �        55
 ���������        55 P        h5{5 �        h5{5 Q        h5{5
 ���������        h5{5 P        �56 R66 P66 R        $6?6 	��?6D6 PD6o6 	��o6q6 Pq6�6 	��        $6D6 � D6p6 Sp6q6 � q6�6 S�6�6 � �6�6 S        �6�6 P        +6D6 � D6p6 Sp6q6 � q6�6 S�6�6 � �6�6 S        2686 1�        2686 �         D6g6 S�6�6 S        ]6g6 S�6�6 S        ]6g6 	���6�6 	���6�6	 s���        86D6 � q6�6 S�6�6 �         <6?6 P        q6�6 S�6�6 �         �6$7 � *7C7 �         �6�6 P        �6�6 S�6�6 � �6(7 S(7)7 � *7C7 S        �6(7 S(7)7 � *7C7 S        77 S*7C7 S        �6�6 P77 	��*7C7 	��        �6�6 R�6�6 r�        �6�6 1�        �6�6 S        P7�7 � �7�7 R        r7t7 P        \7_7 P_7`7 � #        `7�7 � �7�7 R        �7�7 � �7�7 R        �7�7 �        �7�7 P        �7�7 � #@K$"p @K$"-��7�7 � #@K$"� #@K$"-��7�7 r@K$"p @K$"-��7�7 r@K$"q@K$"-��7�7 r@K$"r@K$"-�        �7�7 � �7�7 R        �7�7 	��        �7�7 R        �7�7 Q        �7�7 �{^  �7�7 �{^          	88 P        �78 � 8)8 R)8/8 �         �7	8 	��        �7	8 �         8	8 Q        08i8 � i8q8 R        08o8 �        J8L8 P        58i8 � i8q8 R        C8J8 1�        C8J8 �         G8J8 ��_          �8�8 � �8�8 pd�        �9�9 �         �9�9 S�9�9 � �9�9 S�9�9 � �9�9 S�9�9 �         �9�9 1�        �9�9 S        �9�9 S�9�9 �         �9�9 	���9�9	 s���        �9�9 1�        �9�9 S�9�9 �         :P: � P:T: pd�        :L: �L:T: rd�        �:�: S�:�: �         .;5; 1�        .;3; P3;5; �        P;_; �        T;_; �        T;_; � #        {;�; R�;�; �        {;�; p��;�; � #�        {;~; p        �;�; �        ?<P< SP<Q< P        �<�< S�<�< � �<�< S        �<�< V�<�< V        �<�<  �        �<�< V�<�< V        �<�<  �        �<�< V        �<�< P== P        �<�< S�<�< � �<= S== � =L= S        �<= S== � =L= S        �<= V=L= V        �<G=  �        �<= V=G= V        =G=  �        =G= V        e=|= S=�= S�=�= S        i=x= Qx== �=�= Q�=�= ��=�= Q�=�= �        i=x= Rx=}= V}== �=�= R�=�= V�=�= P�=�= R�=�= V        i=|= S=�= S�=�= S        �=�= P�=�= P        �=> S
>:> S:><> � =>B> S        �=�= V�=> P>
> �
>+> V+><> P        �=> S
>:> S:><> �         
>+> V+><> P        
>:> S:><> �         s?�? u�?�? t�?@ u        �?�? u�?�? t�?@ u        �?�? W�?@ W        �?�? P�?�? uT�?@ uT        �C�C ����C�C P�C�C ���        D
D S
DD uDD t        _DqD RqD�D �        _DyD SyD{D � {D�D S        �D�D ��D�D p �D�D �        �D�D R�D�D �        �D�D S�D�D �         VEXE 0�XEyE P        �F�F 0��F�F P        )HVH SVHXH � XH|H S|H~H �         �H�H 	���H�H V�H�H P�H�H 	���H�H V�H�H P�H I V        �H�H � #,80.�        �H�H � �H I S        �H�H P�H�H P        �H�H P        �H�H P         I*I 0�*I.I P        II RI*I �         I%I P        6I5J 	��>JWJ 	��WJYJ VYJ~J 	��        6IjI � #,80.��I�I s,80.�        XI�I W�I&J W>JFJ WFJMJ PMJ~J W        nIsI PJ&J P        XI�I �z{  �IJ �z{  J&J ��{  >J~J �z{          XInI �{  nI�I ��{  �I&J �{  >J~J ��{          dInI �         dInI 	��        jInI Q        �I�I �z{          �I�I 	��        �I�I S        �I�I s,80.�        �I�I P        �I�I S        UJYJ �z{          �JK 0�KK P#KHK 0�HK�K P�K�K 0�        �J�J P�J�J W�J�J P�K�K W        �J�J P�K�K P        �J�J P        �J#K 
 �HK�K 
 �        �JK R        �J#K �Z~  HK�K �Z~          �J#K �I~  HK�K �I~          �J!K WHK�K W        �J�J P�JK t KK �@        HK�K 0�        HK�K S        HK�K s,80.�        VKbK 0�}K�K 1�        YKwK R�K�K R�K�K s4        YK}K S�K�K S        bKwK 0�        bKwK S        �K�K r q "1��K�K R        �K�K R�K�K s4        �K�K S        �K�K � #,80.��M�M s,80.�        �K�K P�KrM �H�M�M �HN�N �H�NP �H        �K�L 0��L�L W�L�L Q�LAM 0��M�M WNN WN�N 0��N�N W�N�N P�N�N 0�;O�O 0��O�O P�O�O W�OP 0�        �K|L 0�|L�L V�L�L U�L M U M;M 0�;MAM P�M�M UN'N UdNN UN�N V�N�N U�N�N P;O�O 0��O�O U�O P 0� PP UPP 0�        �K|L 0�|L M V MrM 0��M�M VN#N VDNSN PSN�N V�N�N V�N�N 0�;O�O 0��O�O V�O P 0� PP VPP 0�        �K�L � �LrM S�M�M S�M�M � NP S        �N�N S        �N�N R        �N�N P        �N�N s4        �N�N S        �KL PPP P        LL P        9L~L U;O�O U�O P U        9LLL PLL�L W�L�L 1��LM WN�N W;O�O W�OP W        EL|L V;O�O V�O P V        L&L P        ROXO P�O�O P�O P �D        �L�L PM M P        VNhN s� p �        dNnN P        dNnN Q        N'N �\�'N.N U.N1N t 1NAN ��ANSN �\�        N0N q �H"�0NSN U        N5N Q5N6N t 6NAN ��        NSN s� �        NAN R        N;N P;N<N t <NAN ��        NSN s1�        N*N s�         �O�O P        AMrM 	��        AMrM S        AMWM s,80.�        (O;O 0�        (O;O S        PMrM PO:O P        PMrM SO;O S        �M�M U�N�N U        �M�M S�N�N S        �M�M s,80.�        �M�M p u "��M�M U�N�N p u "�        �M�M P�N�N P        �M�M S�N�N S        �M�M 0�        �M�M S        �M�M P        �MN 	��        �MN S        �M�M s,80.�        NN 0�        NN S        �MN P        �MN S         P]P �]PcQ VfQ�Q ��Q�Q V�QR �RR VRR t RvR VyR�R V�R�R ��R�R S�R�R V�R�R S�R�R V         P]P �]P�P U�PQ u p �QeQ UfQ�Q ��Q�Q U�QR �RR UR!R U�R�R ��R�R U         P]P 0�]PbQ SbQfQ PfQ�Q 0��Q�Q S�QR 0�RR SRuR SuRyR PyR�R S�R�R 0��R�R 1��R�R S�R�R 1��R�R S        �P�P w 80.��R�R w 80.�        �P�P P�P�P p81r p8@K$"  �*( ��P�P  � #81r � #8@K$"  �*( ��P�P � #811� #8@K$"  �*( ��R�R  � #81r � #8@K$"  �*( �        ]P�P � �R�R Q�R�R Q        ]P�P �         oP�P R        oP�P P        oP�P � #4        oP�P �         �P�P P�R�R P        �P�P P        �P�P �\p �        �PQ PQ3Q P!R4R P�R�R P        /QfQ 	��        /QfQ �         /QfQ � #,80.�        :QaQ PaQfQ � #4        :QfQ �         \QfQ 0�        \QfQ �         R!R W        RR P        RR VRR t         !R�R 0�        !RyR � yR�R P�R�R �         !RNR � #,80.�yR�R p,80.��R�R � #,80.�        :RNR 0�yR�R 1�        ERRR P�R�R P�R�R q4        ERNR � NRyR Q�R�R Q        NRgR 0�        NRgR �         �R�R p r "1��R�R P        �R�R P�R�R q4        �R�R Q        �Q�Q 	��        �Q�Q �         �Q�Q � #,80.�        �Q�Q P        �Q�Q �         �Q�Q 0�        �Q�Q �         �R�R Q�R�R Q        �R�R 1��R�R 1�        
S)S �         S&S � #@�&S)S R        S&S R&S)S � #        S)S �         ;S_S �         SS_S Q        SS_S R        IS_S S        IS_S �         |S>T S>TAT uATBT tBTcT ScTfT ufTgT tgT�T S        �T�T �         �U�U PV#V PYV^V P        �U�U VV&V V&VYV �Dw �YVcV V        RUbU PsVwV P        ZUbU P        vUyU v p �yU�U P�U�U VV&V V&VdV �Dw �        �U�U W�U�U ��UdV WfVsV W        �U�U P�U�U P�U<V �@<VUV PfVrV P        mUuU P        �U�U R�U�U �X��U&V �X�&V,V V,V-V t -V.V t.V/V t/V2V t2V5V t5V8V t8V9V t9V;V t;VsV �X�        �U�U w p "��U�U P�U�U t �U�U t�U�U t�U�U t�U�U t�U�U t�U�U t        �U�U W�UdV WfVsV W        �U�U �\��U�U P�U�U t �U�U t�U�U t�U�U t�U�U t�U�U �\��U,V �\�,VGV VGVsV �\�        �U�U �v "��U�U P�U�U �v "��UV �v "�VsV ��"�        �U�U ��UsV �        �U�U �L�UsV �L         V,V �\,V;V v          V)V s�\�LVcV V        #V&V �X�&V,V V,V-V t -V.V t.V/V t/V2V t2V5V t5V8V t8V9V t9V;V t;VfV �X�        #V;V R;VfV �D        #VdV W        #V,V �\�,VGV VGVfV �\�        #V)V s        #V,V �\,V;V v         #VfV �L        #V;V P        �V�V P        �V�V S�V�V �         �V�V P        �V�V ss��V�V P        �V�V s�         �V�V s�         �V�V R        �VW 1�WX ��~X;X 1�;X@X ��~        +X;X P        WW P;X?X P        WW P        PWhW S�W�W P�W�W S�W�W P�WX S        PW�W ��~�W�W R�W�W R�W�W ��~        PWhW ��~�kWrW ��~�rW~W Q~W�W ��~��WX ��~�        PWhW UkW�W U�WX UXX �`�        PWhW WkW�W W�WX WXX ��~�        PWhW ��~kW�W ��~�WX ��~        kW~W P        �W�W P        �W�W P        KX{X U{X~X � ~X�X U�X�X �         �X�X P�R��X�X p �R�        �X�X S�X�X �        �X�X s,80.��X�X �#,80.�        �X�X S�X�X �        �X�X S�X�X �        �XqY 1�~Y�Z 1�        Y$Y P        �X5Y S�Y*Z S        �Y*Z S        Z*Z R        Z*Z P        	Z*Z s4        	Z*Z S        IYYY �S�          MYYY S        MYYY 1�        �Y�Y 0��Z�Z 0�        �Y�Y S�Z�Z S        �Y�Y s,80.��Z�Z s,80.�        �Y�Y 0��Z�Z 1�        �Y�Y P�Z�Z P�Z�Z s4        �Y�Y S�Z�Z S        �Z�Z p r "1��Z�Z P        �Z�Z P�Z�Z s4        �Z�Z S        �Y�Y �S�          �Y�Y S        �Y�Y 1�        �Y�Y �S�  �Z�Z �S�          �Y�Y �S�          *Z�Z 0�        *Z�Z S        *Z�Z s,80.�        6ZBZ 0�YZ�Z 1�        9ZYZ PfZ~Z P~Z�Z s4        9ZYZ SfZ�Z S        BZYZ 0�        BZYZ S        tZ~Z p r "1�~Z�Z P        tZ~Z P~Z�Z s4        tZ�Z S        �Z�Z 0��Z[ P[�\ �D        F[�[ V�[�[ Q�[�[ Q�[�[ Vo\x\ V�\�\ V        �Z�Z P        F[�[ S�[�[ ��[i\ Si\o\ �o\�\ S        u[�[ 1��[o\ 0�o\�\ 1��\�\ 0��\�\ 1�        u[�[
 �        �[�[ V�W�"\D\ R�Q�o\z\
 �        z\�\ V�W��\�\ V�W��\�\ R�Q��\�\ R�Q��\�\
 �        �\�\ V�W�        �[�[ P�R�        �[�[ P        �[i\ Si\o\ ��\�\ S        �[\ S        �[\ V        �[\ P        �[\ s4        �[\ S        ]X] SX]\] �\]�] S        �\Y] VY]\] � \]�] V        ]R] S\]�] S        �]�] 1��]b^ 1�b^n^ p 	�.�n^|^ 0�|^�^ 1��^�^ P�^9_ 1�        �]�] 0��]�] V�]�] � #L�]z^ V|^�^ V�^�^ 0��^9_ V        �]�] S�]�] � �]y^ Sy^|^ � |^�^ S�^9_ S        �]�] P        �]�] P        ^#^ P        ^#^ P        3^n^ V        Z^n^ �d�        __ r p �__ R_._ R._4_ W        �^�^ R�^�^ t �^�^ �L        �^�^ s�         �^_ W        �^�^ s2��^�^ R�^4_ s2�        �^�^ P        �^�^ 	��        �^�^ S        �^�^ s,80.�        �^�^ 0�        �^�^ S        �^�^ P        �^�^ S        @_�_ � �_�_ P        @_�_ ��_�_ R        L_U_ q 80.�U_�_ � #,80.��_�_ p,80.�        R_�_ S�_�_ � #,�AH$0.��_�_ S�_�_ p,�AH$0.��_�_ S        X_f_ q �"�f_i_ Qi_�_ � #4�"��_�_ p4�"��_�_ q r "�        X_f_ Qf_�_ � #4�_�_ p4�_�_ Q        X_�_ � �_�_ P        |_�_ q r "1��_�_ R        |_�_ Q        |_�_ �         �_�_ 0�        �_�_ P        �_�_ �         �_�_ � #�        �_�_ �         �_�_ � #�         `` �          `` � #�        `` �         `` � #�        0`5` �         0`5` � #�        @`E` �         @`E` � #�        �`�` 0��`3a VJaqa 0�qa�a 1��a�a 0��a�a 1��a�a 0�        �`2a S2a6a P6aFa SFaHa w\�Ja�a S�a�a u�a�a S�a�a u�a�a w\�        �`2a S2a6a PJa�a S�a�a u�a�a S�a�a u�a�a w\�        �`5a ud�5a6a t`�Ja�a ud�        �`5a ud�5a6a t`�        �`6a 	��        �`a R        �`a r,80.�        a6a 0�        aa R        �`a P        �aQb v�QbSb u#�SbTb t#�Tbb v�        �aPb SPbSb uSbTb tTbb S        �b�b s� ��bc Vcc u#h�cc t#h�cMc V        �bc Scc ucc tcMc S        _c�c v��c�c u#��c�c t#��c�c v�        _c�c S�c�c u�c�c t�c�c S        �c�c s� ��cud Vudwd u#d�wdxd t#d�xd�d V        5dtd Stdwd uwdxd txd�d S        �dGe v�GeIe u#�IeJe t#�Je~e v�~ee u#�e�e V        �dFe SFeIe uIeJe tJe�e S        �dGe v�GeIe u#�IeJe t#�Je~e v�~ee u#�e�e v�        �dGe v�GeIe u#�IeJe t#�Je~e v�~ee u#�e�e v�        �dFe s�FeIe u#�IeJe t#�Je�e s�        Uele v�        Uele S        �e�e s� ��eKf VKfMf u#l�MfNf t#l�Nf�f V        �eqf �	�qfrf t rfvf tvf�f �	�        �eJf SJfMf uMfNf tNf�f S        fNf �	�Rfzf �	�        fJf s�JfMf u#�MfNf t#�Rfzf s�        �f*g 0�*g.g P.gug 0�ugyg P        �f+g S+g.g � .gvg Svgyg �         �f+g S+g.g � .gag S        �fag �        �f-g W-g.g �.gag W        �f+g S+g.g � .gag S        gag 	��        g+g S+g.g � .gag S        g-g w 80.�-g.g �80.�.gag w 80.�        gag 0�        g+g S+g.g � .gag S        g%g P.g2g P2gAg s4        �g�g �        �g�g P�g�g �        �g�g p 8!��g�g �8!�        �g�g ��g�g �        �g�g s��g�g P�g�g s��g�g � #��g�g s��g�g � #�        �g�g �        �g�g S�g�g �         �g�g S�g�g �         �g�g s�g�g P        �g�g P�gLh �        �g�g p @!��gLh �@!�        �gh �0hCh �        �g	h s�	hh Ph#h s�#h'h � #�0h5h s�5h<h � #�        0hCh �        0h5h S5h<h �         5hGh SGhKh �         5h<h s<h?h P        Xhzh ��h�h �        Xheh s�ehjh Pjhh s�h�h � #��h�h s��h�h � #�        �h�h �        �h�h S�h�h �         �h�h S�h�h �         �h�h s�h�h P        �h�h P�hi �        �hi �        �h�h S�h�h �         �hi Sii �         �h�h s�h�h P        ii Pili �        Nici �        NiUi SUi\i �         Uigi Sgiki �         Ui\i s\i_i P        �i�i �        �i�i S�i�i �         �i�i S�i�i �         �i�i s�i�i P        �i�j v��j�j u#��j�j t#��j�j v��j�j u#��j�j t#��j�j v��jk V        �i�j S�j�j u�j�j t�j�j S�j�j u�j�j t�jk S        �i�j v��j�j u#��j�j t#��j�j v��j�j u#��j�j t#��j�j v��jk v�        j�j v��j�j u#��j�j t#��j�j v��j�j u#��j�j t#��j�j v��jk v�        j�j s��j�j u#��j�j t#��j�j s��j�j u#��j�j t#��jk s�        �j�j v�        �j�j S        bj�j u�j�j t�j�j u�j�j t        bj�j u�j�j t�j�j u�j�j t        bj�j S�j�j u�j�j t�j�j S�j�j u�j�j t        �j�j u�j�j t        �j�j u�j�j t        �j�j S�j�j u�j�j t        �j�j 4�        �j�j R        �j�j r        k�k v��k�k u#��k�k t#��k�k v��kl u#�ll t#�l6l v�6lGl V        k�k S�k�k u�k�k t�k�k S�kl ull tlGl S        k�k v��k�k u#��k�k t#��k�k v��kl u#�ll t#�l6l v�6lGl v�        Ak�k v��k�k u#��k�k t#��k�k v��kl u#�ll t#�l6l v�6lGl v�        Ak�k s��k�k u#��k�k t#��k�k s��kl u#�ll t#�lGl s�        l$l v�        l$l S        �k�k u�k�k t�kl ull t        �k�k u�k�k t�kl ull t        �k�k S�k�k u�k�k t�k�k S�kl ull t        �k�k W�k�k u#��k�k t#��k l W ll u#�ll t#�        �kl ull t        �kl ull t        �k�k S�kl ull t        �kl 4�        �k�k R        �k�k r        \l_l s� �_l3m V3m5m u#l�5m6m t#l�6m_m V_mam u#l�ambm t#l�bm�m V        �l�m �	��m�m t �m�m t�m�m �	�        �l2m S2m5m u5m6m t6m^m S^mam uambm tbm�m S        �lbm 0�fm�m 0�        �lbm �	�fm�m �	�        �l2m s�2m5m u#�5m6m t#�6m^m s�^mam u#�ambm t#�fm�m s�        m5m u5m6m t6mam uambm t        m5m u5m6m t6mam uambm t        m2m S2m5m u5m6m t6m^m S^mam uambm t        6mam uambm t        6mam uambm t        6m^m S^mam uambm t        Jmbm 4�        JmVm R        JmQm r        �m�m s� ��m�n V�n�n u#l��n�n t#l��n�n V�n�n u#l��n�n t#l��no V        n�n �	��n�n t �n�n t�no �	�        n�n S�n�n u�n�n t�n�n S�n�n u�n�n t�no S        %n�n 0��n�n 0�        %n�n �	��n�n �	�        %n�n s��n�n u#��n�n t#��n�n s��n�n u#��n�n t#��n�n s�        in�n u�n�n t�n�n u�n�n t        in�n u�n�n t�n�n u�n�n t        in�n S�n�n u�n�n t�n�n S�n�n u�n�n t        in�n W�n�n u#��n�n t#��n�n W�n�n u#��n�n t#�        �n�n u�n�n t        �n�n u�n�n t        �n�n S�n�n u�n�n t        �n�n 4�        �n�n R        �n�n r        o�o v��o�o u#��o�o t#��o�o v��o�o u#��o�o t#��o�o v�        o�o S�o�o u�o�o t�o�o S�o�o u�o�o t�o�o S        do�o u�o�o t�o�o u�o�o t        do�o u�o�o t�o�o u�o�o t        do�o S�o�o u�o�o t�o�o S�o�o u�o�o t        do�o @�        �o�o u�o�o t        �o�o u�o�o t        �o�o S�o�o u�o�o t        �o�o 4�        �o�o R        �o�o r        �otp v�tpvp u#�vpwp t#�wp�p v��p�p u#��p�p t#��p�p v�        �osp Sspvp uvpwp twp�p S�p�p u�p�p t�p�p S        Dpvp uvpwp twp�p u�p�p t        Dpvp uvpwp twp�p u�p�p t        Dpsp Sspvp uvpwp twp�p S�p�p u�p�p t        Dp�p @�        Dpvp u@!�vpwp t@!�wp�p u@!��p�p t@!�        Dpup Wupvp u#�vpwp t#�wp�p W�p�p u#��p�p t#�        wp�p u�p�p t        wp�p u�p�p t        wp�p S�p�p u�p�p t        �p�p 4�        �p�p R        �p�p r        �p]q v�]q_q u#�_q`q t#�`qq v�q�q u#��q�q t#��q�q v�        �p\q S\q_q u_q`q t`q~q S~q�q u�q�q t�q�q S        /q_q u_q`q t`q�q u�q�q t        /q_q u_q`q t`q�q u�q�q t        /q\q S\q_q u_q`q t`q~q S~q�q u�q�q t        /q�q 8�        `q�q u�q�q t        `q�q u�q�q t        `q~q S~q�q u�q�q t        jq�q 4�        jqvq R        jqqq r        �q?r v�?rAr u#�ArBr t#�Bror v�orqr u#�qrrr t#�rr�r v�        �q>r S>rAr uArBr tBrnr Snrqr uqrrr trr�r S        rAr uArBr tBrqr uqrrr t        rAr uArBr tBrqr uqrrr t        r>r S>rAr uArBr tBrnr Snrqr uqrrr t        rrr 8�        rAr u8!�ArBr t8!�Brqr u8!�qrrr t8!�        r@r W@rAr u#�ArBr t#�Brpr Wprqr u#�qrrr t#�        Brqr uqrrr t        Brqr uqrrr t        Brnr Snrqr uqrrr t        Zrrr 4�        Zrfr R        Zrar r        �r�r s� ��ras Vascs u#d�csds t#d�ds�s V�s�s u#d��s�s t#d��s�s V        �r`s S`scs ucsds tds�s S�s�s u�s�s t�s�s S        3scs ucsds tds�s u�s�s t        3scs ucsds tds�s u�s�s t        3s`s S`scs ucsds tds�s S�s�s u�s�s t        3s�s @�        ds�s u�s�s t        ds�s u�s�s t        ds�s S�s�s u�s�s t        zs�s 4�        zs�s R        zs�s r        �s�s s� ��s�t V�t�t u#d��t�t t#d��t�t V�t�t u#d��t�t t#d��t�t V        t�t S�t�t u�t�t t�t�t S�t�t u�t�t t�t�t S        St�t u�t�t t�t�t u�t�t t        St�t u�t�t t�t�t u�t�t t        St�t S�t�t u�t�t t�t�t S�t�t u�t�t t        St�t @�        St�t u@!��t�t t@!��t�t u@!��t�t t@!�        St�t W�t�t u#��t�t t#��t�t W�t�t u#��t�t t#�        �t�t u�t�t t        �t�t u�t�t t        �t�t S�t�t u�t�t t        �t�t 4�        �t�t R        �t�t r        �t�t s� ��t�u V�u�u u#h��u�u t#h��u�u V�u�u u#h��u�u t#h��u v V        5u�u S�u�u u�u�u t�u�u S�u�u u�u�u t�u v S        zu�u u�u�u t�u�u u�u�u t        zu�u u�u�u t�u�u u�u�u t        zu�u S�u�u u�u�u t�u�u S�u�u u�u�u t        zu�u 8�        �u�u u�u�u t        �u�u u�u�u t        �u�u S�u�u u�u�u t        �u�u 4�        �u�u R        �u�u r        vv s� �v�v V�v�v u#h��v�v t#h��v�v V�v�v u#h��v�v t#h��v w V        Uv�v S�v�v u�v�v t�v�v S�v�v u�v�v t�v w S        �v�v u�v�v t�v�v u�v�v t        �v�v u�v�v t�v�v u�v�v t        �v�v S�v�v u�v�v t�v�v S�v�v u�v�v t        �v�v 8�        �v�v u8!��v�v t8!��v�v u8!��v�v t8!�        �v�v W�v�v u#��v�v t#��v�v W�v�v u#��v�v t#�        �v�v u�v�v t        �v�v u�v�v t        �v�v S�v�v u�v�v t        �v�v 4�        �v�v R        �v�v r        Hw\w S        HwOw s        �w�w S        �w�w s        �w�w S        �w�w s        �wx Sxx �         �wx Sxx �         :x=x s�=xIx PIxyx s�yx{x � #�        Uxyx s�yx{x � #�        gxzx v�zx{x �#�        gxyx Syx{x �         �x�x s��x�x P�x�x s��x�x � #�        �x�x s��x�x � #�        �x�x v��x�x �#�        �x�x S�x�x �         �xy Pyy s�y/y � #�/y3y s��3y7y � `�        yy s�y/y � #�/y3y s��3y7y � `�        hyty Pty�y s��y�y � #��y�y s���y�y � `�        �y�y s��y�y � #��y�y s���y�y � `�        �y�y s��y�y P�yCz s�CzEz � #�        �yCz s�CzEz � #�        zDz v�DzEz �#�        zCz SCzEz �         !zDz v�DzEz �#�        !zCz s�CzEz � #�        1zDz v�DzEz �#�        1zCz SCzEz �         Xz�z S�z�z �         hztz Ptz�z s��z�z � #�        �z�z s��z�z � #�        �z�z s� ��z�z P�z�z s� ��z�z � #d�        �z,{ S,{0{ �         �z�z P�z,{ s�,{0{ � #�         {,{ s�,{0{ � #�        {{ s� �{#{ P#{,{ s� �,{0{ � #h�        o{{{ P{{�{ s��{�{ � #��{�{ s���{�{ � `�        �{�{ s��{�{ � #��{�{ s���{�{ � `�        �{3| S3|7| �         �{�{ P�{3| s�3|7| � #�        |3| s�3|7| � #�        || s� �|*| P*|3| s� �3|7| � #l�        p}�} � �}�} R�}�} R        p}�} ��}�} Q�}�} Q        p}�} ��}�} P�}�} P�}�} �        �}�} ��}�} P        �}�} ��}�} Q        �}�} � �}�} R        �}�} � �}�} R�}�} R        �}�} ��}�} Q�}�} Q        �}�} ��}�} P�}�} P�}�} �        �}�} ��}�} P        �}�} ��}�} Q        �}�} � �}�} R        �}~ � ~~ Q~#~ Q        �}~ �~~ R~#~ R        �}~ �~#~ �        ~~ P        ~~ �~~ R        ~~ � ~~ Q        0~O~ � O~S~ QT~f~ Q        0~4~ �4~S~ RT~f~ R        <~>~ P>~G~ �T~f~ �        <~S~ �T~f~ �        <~O~ � O~S~ QT~f~ Q        >~S~ PT~c~ Pc~f~ ���        >~S~ �T~f~ �        >~O~ � O~S~ QT~f~ Q        C~S~ P        C~S~ �        C~O~ � O~S~ Q        p~�~ � �~�~ Q�~�~ Q        p~t~ �t~�~ R�~�~ R        |~~~ P~~�~ ��~�~ �        |~�~ ��~�~ �        |~�~ � �~�~ Q�~�~ Q        ~~�~ P�~�~ P�~�~ ���        ~~�~ ��~�~ �        ~~�~ � �~�~ Q�~�~ Q        �~�~ P        �~�~ �        �~�~ � �~�~ Q        �~�~ � �~�~ Q�~�~ Q        �~�~ ��~�~ R�~�~ R        �~�~ ��~�~ �        �~�~ P�~�~ P�~�~ �r �        �~�~ ��~�~ R�~�~ R        �~�~ � �~�~ Q�~�~ Q        �~�~ P        �~�~ ��~�~ R        �~�~ � �~�~ Q        �~ �  Q& Q        �~ � R& R        �~ �& �        �~ P# P#& �r �        �~ � R& R        �~ �  Q& Q         P         � R         �  Q        08 � ��89 P        PZ F�Z[ �         lr F�rs �        ��	 r rt"���� R�        �� ���� R�        ��	 r rt"���"� R�        8�<� ��<�?� R�        �� pt1��� r�        ��� �P�a� �        ��� P�P� �P�`� P`�a� �        	�(� R(�3� �3�G� RG�P� �        	�� P�P� �        	�P� �         	�� s p @K$"r @K$"+��� qtp @K$"r @K$"+��(� qt�@K$"r @K$"+�3�G� qt�@K$"r @K$"+�G�I� qt�@K$"�@K$"+�        �,� S3�O� SO�P� P        �(� P3�C� PC�P� q �"�        �,� �3�P� �        �,� S        �(� P        �,� �        C�P� �        p��� � ���� S        p��� ����� Q        u��� � ���� S        ���� �        ���� pt�        ���� P        ���� �         ���� R        ���� �         �F� �N��� ����� P���� Q��ʂ �TʂՂ PՂڂ q�ڂ� Q        '�N� � N�W� PW�� �         ��ʂ �1�ڂ� �1�        ��ʂ �#�ڂ� �#�        ��ʂ Vڂ� V        �4� S4�5� �        C�]� 	��]�`� S`�c� Pc��� 	������ S���� P        c�u� q ��u��� Q        c�z� v �"�z��� R���� v �"�        ��ۃ �ۃ� S�� P�� S�� P�� s�        ݃� V�� ��� V�� �        ݃� U�� ��� U�� �        ݃� w s "���� P��� w s "��� w p "��� w s "�        H�d� Sd�e� �        p��� ����� S���� �        ���� P���� P        ��Ԅ �Ԅ� S�&� S&�*� P        ؄� � �*� �         ��� w s "��� w s "1��&� w s "�&�(� w p "�        ��� V�'� V'�*� �        ��� ��*� �        X�t� St�u� �        ���� ����� P        Å̅ S̅΅ vt1�΅Յ SՅم Pم�� S���� P        ���� � ��΅ P΅�� �         ΅�� v s "����� v p "�        ΅�� W���� �        ΅�� U���� �        (�D� SD�E� �        P�Y� �Y�]� P        `�o� �o��� V���� P��ʆ V        o�|� P|�͆ �         ���� s v "����� s v "1����� s v "�        ���� W���� �        ���� U���� �        ��� S�� �         �D� �D�a� P        ���� S���� vt1����� S���� P��Շ SՇ� P�� s�        ��Շ v s "�Շև v p "�ه� v s "�        ��؇ U؇ه �ه� U�� �        ��ׇ Wׇه �ه� W�� �        �4� S4�5� �        @�Z� �Z��� S���� �        c�l� Pl�n� r�n�u� Pu�y� Ry��� P���� R        ���� S���� pt        �� V        ���� R        ���� P        Ј� ��*� R*�+� �        Ј� ��� S��+ � <��� <�@K$"�@K$",( ��*� Q*�+� �        ��� V        �� P        ߈� ��*� R*�+� �        �� �        �� �        �� �         �� s �@K$"�@K$"+��� pt�@K$"�@K$"+��� � <�@K$"�@K$"+�        �� �        ��� Q        ��� p �"��� P        0�d� �d��� S���� �        0�o� �o��� R���� �\���� �        ���� P        C��� Q���� ����� Q���� ����� Q���� �        C�T� RT��� � ���� R���� �         P��� �	����� �	�        P�� V��� ����� V        P��� ����� �        ]�t� Pt��� �        ]��� Q���� �        ]��� �         ]�_� s q @K$"p @K$"+�_�t� wtq @K$"p @K$"+�t��� wtq @K$"�@K$"+����� wt�@K$"�@K$"+�        d��� �        d�� V��� �        d��� �        d�f� r v @K$"�@K$"+�f�� utv @K$"�@K$"+���� ut�@K$"�@K$"+�        o�� u v "���� V���� u �"�        o��� w q "����� Q���� w �"�        ԉ� S        ߉� P��� V        ԉ�� U���� �        ߉�� U���� �        ߉�� W         �#� �#�A� SY�j� �        4�<� P<�W� W        Q�Y� P        �V� VV�Y� �Y�j� V        �Y� � Y�i� Ri�j� �         �Y� � Y�i� Ri�j� �         �.� P.�Y� �        �V� VV�Y� �        �Y� �         �� s v @K$"p @K$"+��.� utv @K$"p @K$"+�        #�Y� �        4�Y� �        4�:� u v "�:�K� RK�V� u v "�V�X� u �"�        p��� ����� S����) � <r �� <r @K$"�@K$",( ���ʊ �        ���� P        }��� R���� ���Ɋ RɊʊ �        ���� Q���� �        ���� R���� �        ���� �         ���� s r @K$"q @K$"+����� ptr @K$"q @K$"+����� ptr @K$"�@K$"+����� � <r @K$"�@K$"+�        ���� �        ���� p r "����� P        p��� � ���� S���� s�`���؋ S؋ً pً� �         ��ً 
 �        ��ً @�        ���� s����� s�`�����! � �1$� @K$"�1$@K$"*( #���ɋ R        ���� R���� s�`�����! � �1$� @K$"�1$@K$"*( #�        ʋً P        ���� 
 r 
������ 
 s�`
������) 
 � �1$� @K$"�1$@K$"*( #
��        ��ً 0�        ��ɋ R        ͋ً P        �?� �I�p� �        �,� U,�3� P3�7� UI�W� U        �?� SI�p� S        �&� P&�?� WI�R� PR�p� W        "�,� U,�3� P3�7� UI�W� U        "�?� SI�p� S        "�?� VI�p� V        $�,� U,�3� P3�7� U        $�7� S        $�7� V        I�W� ��Q          I�W� V        7�?� SW�p� S        7�?� WW�p� W        ���� ����� P        ��Č	 � ##�        Ќ�� P��� �P�        Ќ�� R��� �R�        Ќ�� p���� �P#�        ׌�� Q��� s�        #�2� Q        M�t� �o�t�z� Pz��� �o�        M�U� RZ�z� R        Z�t� �o�t�z� Pz��� �o�        Z�z� R        Z�z� r�        c�z� Qz��� s�        ��+� U,��� U��C� U        ��� V,��� V��#� V        ͍Ӎ PӍ� Q�� P��� Qَ� Q��� �L        ύ� � َ�� �         ۍ� Wَ�� W        ۍ� P�� � َ� P        ۍ� Rَ� R��� �H        �� R        ��� W        �� P        �� R��� �H        ۍ� Qَ� Q��� �L        ��� � �C� �         �� S�� �_��C� S        �� Q�:� Q        �:� Q        �:� q�        �� �H        �� �         F�V� V��� V        F�R� PR�T� � �"�"���
� P        F�V� Q��
� Q        R�V� Q        ��� V        ��
� P        ��
� Q        |��� V��َ V        |��� P���� � �"�"���ʎ P        |��� S��Ԏ S        ���� S        ��َ V        ��ʎ P        ��Ԏ S        �+� U���� U        �$� st����� st�        ���� U        ���� s u "�        y��� pt�        ���� � <����� rt�        ͏� S��� �        �� V��� P        ��� S� � �        �� V� � P        -�O� SO�S� �        D�P� VP�S� P        ѐ� S        ��#� � #�0� V        �#� �         =�_� S_�c� �        T�W�	 r rt"��W�c� R�        T�`� V`�c� P        w��� P���� �         ��đ Vđő �ő֑ V        ���� Q��ő �őՑ QՑ֑ �        ��ő � ő֑ S        ���� p q @K$"v @K$"+�őՑ p q @K$"v @K$"+�        ��ő � ő֑ S        ���� Q��ő �őՑ QՑ֑ �        ��ő � ő֑ S        ��� ��� S        �� S        ��� pt��� �<�         �(� �(�X� R        0�2� q ��2�X� QX�x� ���        L�u� S        _�o� rt�o�x� �<�        ��ޒ Sޒ� ���� S���� ���� S        ���� P���� ���
� P
�� �        ��ߒ Vߒ� � ��� V���� � ��� V        ��ؒ ���� �        ��͒ U͒Ԓ PԒؒ U��� U        ��ؒ S��� S���� �        ���� W��ؒ ���� �        ��ؒ V��� V���� �         ��͒ U͒Ԓ PԒؒ U��� U        ��ؒ S��� S���� �        ��ؒ W��� W        Œ͒ U͒Ԓ PԒؒ U        Œؒ S        Œؒ W        ��� �f          ��� W        �-� P-�2� �         M�c� Sc�d� P        ���� P���� ����� P���� �        ���� R���� � ���� R���� �         ��ϓ �ϓԓ S        ԓ� S        ��� pt����� �<�         �:� � N�_� �          �B� �N�_� �         �>� �N�_� �         �6� �N�_� �         �2� �N�_� �        �I� UN�_� U        �M� RN�^� R^�_� �        �F� SF�M� � N�_� S        !�I� q r @K$"u @K$"+�N�^� q r @K$"u @K$"+�        *�M� RN�^� R^�_� �        *�F� SF�M� � N�_� S        `�i� �i�}� P        `�q� �q�u� Ru��� �        ���� ����� P        ���� R���� �         ��� � �� �        ��� � �� S�� �        ��� � �� �        ��� � �� �        ��� �  �� W�� �         ��� � �� S�� �        ��� � �� �        ��� V �� V        ��� �        ��� �        ��� V        �� V        �P� � P�~� S~��� � ��ƕ S        �P� �P�n� Pn��� ����� P���� ����� P���� ���ŕ Pŕƕ �        �P� �P�ƕ V        �L� � L�M� SM�P� � P�~� S~��� P��ƕ S        *�L� �L�N� VN�P� �P�ƕ V        *�H� QP�Y� QY�h� rt���� rt���� rt��ŕ Q        *�L� � L�M� SM�P� � P�~� S~��� P��ƕ S        0�P� �P�n� Pn��� ����� P���� ����� P���� �        0�L� � L�M� SM�P� � P�~� S~��� P���� S        [�n� Q���� Q���� Q        _�t� V        _�n� Pn�t� �        _�n� R        d�t� V        d�n� Pn�t� �        d�n� R        t��� V        t��� rt�        ~��� V        ~��� rt�        ���� r v "�        ���� V        ���� P���� �        ���� R        ���� V        ���� P���� �        ���� R        ���� R        �� � �%� V%�*� � +�<� V        �#� �+�<� �        �� �+�;� P;�<� �        �+� �+�<� S        �+� �+�<� S        �� �+�;� P;�<� �        �#� �+�<� �        �� q �@K$"�@K$"+�+�;� q p @K$"s @K$"+�        �� �+�;� P;�<� �        �#� �+�<� �        H�`� S`�a� �        ���� S���� �        ���� � �#� �#�;� RI�f� R��� R��� R�!� �        ���� W �%� W%�x� ���� ����� ���� ��!� W        ���� � ���� S �E� SE�I� � I��� S���� P��!� S        ���� � ���� S �E� SE�I� � I��� S���� P��!� S        Ԗ� 	��!� 	�        Ԗ�� V �F� VF�I� �I�j� Vj�x� ���� V��ŗ Vŗ� ��� V�!� V        Ԗ� 0��!� 0�        Ԗ�� � ���� S �E� SE�I� � I��� S���� P��� S�!� S        ��� R���� � �� R�x� ���� ����� ���� �        ��� � ���� S �E� SE�I� � I��� S���� P��� S        �� R�H� UI�V� U��� U��ŗ U        %�G� WI�l� W��� W��ŗ W�� W        �E� SE�I� � I��� S���� P��� S        ,�F� VF�I� ����� V        ,�;� R���� R        ,�G� W���� W        1�F� VF�I� �        1�;� R        1�G� W        ���� W        X�� Uŗ� U        X�f� R��� R        X�l� W�� W        d�f� W        �� U        ��� R        �� W        n�v� Pv�x� �u �ŗڗ Pڗ� �u �        l�� Vŗ� V        l�� Wŗ� W        v�� W        ŗڗ Pڗ� �u �        ŗ� V        ŗ� W        ��� V��ŗ V        ��� P���� r v "����� P        ��� W��ŗ W        ���� W        ��ŗ V        ���� P        ��ŗ W        0�8� �8�:� P        P��� � ���� �         P��� ����� �        P��� ����� �        P��� ����� �        k��� U���� ����� U        k�� P��� ����� P���� �        k�r� Rr��� ����� �        p�� q p @K$"u @K$"+���� q �@K$"u @K$"+����� q p @K$"u @K$"+�        y�� P��� ����� P���� �        y��� ����� �        ��Ԙ SԘ՘ �        �� pt�� t ��� �h        �"� � "�2� Q2�3� �         �� R"�2� R        �"� � "�2� Q2�3� �         @�O� � O�W� PW�X� �         K�O� � T�W� PW�X� �         O�W� p�W�X� � #�        g�n�	 �� "�        ���� P���� V���� pt���� V�� pt�        ���� R��љ R        ���� � #����� P���� � #���ә s�        ���� P���� W��ę Pęә W        ���� R        ���� � #����� P���� � #�        ���� P���� W        ęә W        ���� V��ә V        ���� � ��ә S        ���� Rљ� R        ���� V���� pt�ϙ� V�� pt�        ә� V�� pt�        ܙ� v r "#��� p r "�        �	� �	�� p @K$"q @K$"+( ��!� �@K$"q @K$"+( �<�I� �        ��8� S8�<� � <�t� S        "�2� PI�j� Pj�t� �L        �4� SI�t� S        	�4� SI�t� S        "�4� SI�t� S        *�2� QI�j� Q        I�j� Q        I�j� q�        2�4� P        2�4� S        ���� R���� u���� t���� u�� t        ߚ.� V.�1� �1�p� V        �'� U1�p� U        �'� S1�p� S        �'� WH�p� W        �� QH�W� Q        �� PH�W� P        �� W        �� Q        �� P        S�W� P        �'� SW�p� S         �'� UW�p� U         �'� pt�W�p� pt�        ���� �0�A� �        ���� W���� ���A� W        ���� Q��0� �0�@� Q@�A� �        ���� P��0� �        ���� W���� ���0� W        ���� Q��0� �        ���� s w @K$"p @K$"+����� rtw @K$"p @K$"+����� rtw @K$"�@K$"+���� rtw @K$"�@K$"+�        ���� U��0� U        ���� V��0� V        ؛�� S�0� S        ؛� R�� R        ؛� P�� P        ݛ� S        ݛ� R        ݛ� P        �� P        ��� V�0� V        ��� U�0� U        ��� pt��0� pt�        �0� U        �0� pt�        *�0� p u "�        g��� S��� S        g��� W��� W��� ���� W        g��� V��� V        ~��� U��� U        g��� H	���� H	�        g��� 0���� 0�        ���� Wǜ͜ W��� W��� �        ���� Vǜ͜ V���� V        ��� W        ��� V        ���� S͜�� S��� S        ���� W͜�� W��� W        ���� R͜ڜ R        ���� R        ͜�� S        ͜�� W        ͜ڜ R        ���� V��� V        ���� U��� U        ���� pt���� pt�        ��� U        ��� pt�        
�� p u "�        8�P� SP�Q� �        x��� S���� �        ��� W��� Q���� W�&� W@�M� W        ��� V�M� V        ��� S�M� S        ʝ� U�@� U        ��� H	��M� H	�        ��� 0��M� 0�        �� W��� Q���� W�&� W        �� V�@� V        ��� P�&� P        �� W��� Q���� W        ��� V        ��� P        �&� ��          �&� P        ��� S&�@� S        ��� U&�@� U        ��� pt�&�@� pt�        &�@� U        &�@� pt�        :�@� p u "�        P��� � ��Ǟ �         P��� ���Ǟ �        P��� ���Ǟ �        X��� Q���� � ���� Q��ƞ QƞǞ �         j��� P���� ����� P���� ���ƞ PƞǞ �        j��� R���� q <���� R��ƞ R        j��� Q���� � ���� Q��ƞ QƞǞ �         ���� 	��        ���� P���� �        ���� Q���� �         ���� 0�        �1� V3�P� V        ��!� � !�0� S0�3� � 3�O� SO�R� �         !�J� ��          !�(� p r "�        &�0� S0�3� � 3�O� SO�R� �         (�1� V3�P� V        3�P� V        J�P� p v "�        k��� W��ğ Q        g��� � ���� S���� � ���� S��ğ �         s��� V�� V        k��� � ���� S���� � ���� S��ğ �         ���� �          ���� r p "�        ���� S���� P���� S��ğ �         ���� V�� V        ���� pt����� s <����� p <����� pt�        �� V        ���� pt�        ���� p v "�        П� � �� P�� P        П�� ���� Q�� Q        П�� ��� �        ԟ� � �� P�� P        ߟ� � �� P        �� �         ��� �        �� �        �� P        /�Y� �o�Y�_� P_�x� �o�        /�_� Qm�x� Q        3�E� Qm�x� Q        E�Y� �o�Y�_� P_�m� �o�        E�_� Q        ;�E� � c�m� �         ���� R��� �        ���� V���� � ��� V        ���� �o���Ԡ �o�Ԡڠ Pڠ� �o��� P�� �o�        ���� Q�� Q��� st���� Q        ���� Q��� Q        �� �o��� P��� �o�        �� Q��� st�        ���� R���� ���� �        ���� V��� V        ���� �o���Ԡ �o�Ԡڠ Pڠ� �o�        ���� R��ڠ R        ��Ԡ �o�Ԡڠ Pڠ� �o�        ��ڠ R        ��� 	��        ��ڠ r�        àڠ Qڠ� w�        ���� V        ,�r� Wr�s� us�v� tv��� W        8�s� us�v� tv��� u        8�B� F�B�L� s L��� F�        B�q� Vq�s� us�v� tv�x� Vx��� u        x��� u        }��� ug����� R���� ug�        }��� P        ��� u�� t�
� u        ���� F���¡ s ¡� F�        ��� W�� u�� t�� W        �
� u        ��� ug��� R�� ug�        ��� P        D�N� uw�N�R� RR�\� uw�        D�R� P        `��� � ��ܢ Vܢߢ � ߢ� V        `�o� �o�x� PȢۢ P        ���� P���� S���� �v ����� �� ���Ȣ Sߢ� S        ���� P���� W���� ut����� pt���â PâȢ Wߢ� W        s�Ȣ ��ߢ� ��        s��� V����� � ���Ȣ V�ߢ� V�        s�Ȣ �y�  ߢ� �y�          s�Ȣ �p�  ߢ� �p�          ��Ȣ ��ߢ� ��        ���� V����� � ���Ȣ V�ߢ� V�        ���� U���� P��Ȣ Uߢ� U        ��Ȣ �ߢ� �        ���� V���� � ��Ȣ Vߢ� V        ���� S���� �v ����� �� ���Ȣ Sߢ� S        ���� S        ���� V        ���� U        âȢ U        ���� S���� �v ����� �� �ߢ� S        ���� W���� ut����� pt�ߢ� W        �h� ���� �        �%� P%�h� ���� �        �]� V]�`� � `�h� V��� V        -�2� P2�\� S\�]� �v �]�`� �� �`�h� S��� S        ;�J� PJ�^� W^�_� ut�_�`� pt�`�c� Pc�h� W��� W        >�h� ���� �        >�]� V]�`� � `�h� V��� V        >�_� U_�`� P`�h� U��� U        >�\� S\�]� �v �]�`� �� �`�h� S��� S        @�N� S        @�N� V        @�N� U        c�h� U        N�\� S\�]� �v �]�`� �� ���� S        N�^� W^�_� ut�_�`� pt���� W        ��ң Vңӣ �ӣ� V        ���� R��ӣ �ӣ� R�� �        ���� s r @K$"v @K$"+����� s �@K$"v @K$"+���ƣ qt�@K$"v @K$"+�ӣ� s r @K$"v @K$"+��� s �@K$"v @K$"+�        ���� R��ӣ �ӣ� R�� �        ���� �o���ѣ Sѣӣ �o�        ��ƣ P        ���� q r "���ƣ R        ǣӣ P        ǣӣ �          �� R�� ��.� R.�/� �         �� Q�� ��.� Q.�/� �        A�H� PH��� �        C�q� Vq�r� �r��� V        C�Y� RY�r� �r��� R���� �        C�H� PH��� �        F�Y� s r @K$"v @K$"+�Y�p� s �@K$"v @K$"+�r��� s r @K$"v @K$"+����� s �@K$"v @K$"+�        S�Y� RY�r� �r��� R���� �        W�r� �        W�e� P        W�Y� q r "�Y�e� R        f�r� �        f�r� P        f�r� �         ��� ��0� �        ��Ť PŤ� ��0� �        ���� V�� � �  �� V�0� V        ͤҤ PҤ�� S���� �v ��� � �� � �� S�0� S        ۤ� P��� W���� ut��� � pt� �� P�� W�0� W        ޤ� ��0� �        ޤ�� V�� � �  �� V�0� V        ޤ�� U�� � P �� U�0� U        ޤ�� S���� �v ��� � �� � �� S�0� S        �� S        �� V        �� U        �� U        ��� S���� �v ��� � �� ��0� S        ��� W���� ut��� � pt��0� W        7�C� p �"�C�I� RI�T� ��"�        7�I� PI�T� �        `��� �̦ݦ �        ץ�� uv "@K$"p w "@K$",����� uv "@K$"uw "@K$",�M�X� uv "@K$"p w "@K$",�X�^� uv "@K$"uw "@K$",����� uv "@K$"p w "@K$",����� uv "@K$"uw "@K$",�        o�¥ W¥å uåĥ tĥr� Wr��� u���� t���� u���� t���� W        c�å uåĥ tĥ�� u���� t���� u���� t���� u        o�å uåĥ tĥ�� u���� t���� u���� t���� u        �å uåĥ tĥ�� u���� t���� u���� t��̦ uݦ�� u        �¥ W¥å uåĥ tĥr� Wr��� u���� t���� u���� t��̦ Wݦ�� W        �å uåĥ tĥ�� u���� t���� u���� t��̦ uݦ�� u        ��� q w @K$"u@K$"+����� ptw @K$"u@K$"+�ĥ�� ptw @K$"u@K$"+����� u<w @K$"u@K$"+�M�X� ptw @K$"u@K$"+�X�Y� u<w @K$"u@K$"+����� ptw @K$"u@K$"+����� u<w @K$"u@K$"+���˦ q w @K$"u@K$"+�        ��̦ 	�ݦ�� 	�        ���� V��å uåĥ tĥ+� V+�M� uM��� V���� u���� t���� V���� u���� t��̦ Vݦ�� V        ���� Sĥ(� SM��� S���� S��̦ Sݦߦ S        ��å uåĥ tĥ�� u���� t���� u���� t��̦ uݦ�� u        ��å uåĥ tĥ�� u���� t���� u���� t���� uݦ�� u        ��å uåĥ tĥ�� u���� t���� u���� t���� uݦ�� u        �M� ud�        �8� uc�8�A� PA�M� uc�        �A� Q        %�8� uc�8�A� PA�M� uc�        %�A� Q        %�M� 	��        %�A� q�        (�M� S        �� uc��� R��� uc�        �� P        X��� uT���� tP���� uT���� tP���� up ����� R���� P        c��� u���� t���� u���� t        r��� V���� u���� t���� V���� u���� t        r��� Q        r��� W���� W        z��� W        ���� V���� u���� t        ���� Q        ���� W        0�o� � ���� �         0�k� ����� �        0�g� ����� �        0�w� ����� �        0�s� ����� �        K�c� Pc�s� ����� P���� �        K�R� RR�w� ����� �        P�c� q p @K$"�@K$"+�c�s� q �@K$"�@K$"+����� q p @K$"�@K$"+�        ]�c� Pc�s� ����� P���� �        ]�w� ����� �        ��ǧ Sǧȧ �        Чԧ �ԧ� P        ��� ���� P        ��� R�� �        �� rt�� t �� �\        �	� R	�� t �� �X        �� Q�� �          �/� �/�E� S        8�@� P@�K� �`        `�d� �d�|� P        `�l� �        ���� ����� P        ���� �        ��Ĩ �ĨԨ P        ̨Ψ R�ΨҨ ��        ̨ب ��        �� ���� P        �� ��� R        �� ��,� P        �� �� � R        Q�_� S        _�k� P        _�v� Sv�w� �        ���� ����� P���        ���� ��"����� R���� ��"�        0�A� PA�F� �P�F�N� PN�T� �P�        0�A� RA�F� �R�F�N� RN�T� �R�        0�A� p�A�F� �P#�F�N� p�N�T� �P#�        7�A� QA�E� s�F�F� QF�T� s�        j��� P        ���� P        ʪ� P        ��� P        S�z� V        V�z� us�        V�]� Pp�w� P        ���� us����� R���� us�        ���� P        �
� V        �
� us�        �� P �� P        %�/� us�/�3� R3�6� us�        %�3� P        s��� V        v��� us�        v�}� P���� P        ���� us���ì RìƬ us�        ��ì P        �*� V        �*� us�        �� P �'� P        E�O� us�O�S� RS�V� us�        E�S� P        ���� V        ���� us�        ���� P���� P        խ߭ us�߭� R�� us�        խ� P        �&� R         �@� V@�A� t A�E� tE�G� t	��G�H� t	��H�I� t	��I�J� t	��J�U� t	��U�b� t	��b�g� t	��g�l� t	��l�m� t	��m�r� t	��r�|� t	��|�~� t	������ t	��         �&� P&��� ��        U�|� V        X�u� �k�u�y� Ry�|� �k�        X�_� Pr�y� P        ���� �k����� R���� �k�        ���� P        �
� V        �
� us�        �� P �� P        %�/� us�/�3� R3�6� us�        %�3� P        s��� V        v��� us�        v�}� P���� P        ���� us���ï RïƯ us�        ��ï P        �*� V        �*� us�        �� P �'� P        E�O� us�O�S� RS�V� us�        E�S� P        ���� V        ���� us�        ���� P���� P        հ߰ us�߰� R�� us�        հ� P        �J� V        &�J� us�        &�-� P@�G� P        |�~� W�P�~�ѱ W�V�ѱ� W���� W�V���� W��        ��ϱ ud�        ��ϱ uc�        ���� Pű̱ P        ��� uc����� R���� uc�        ��� P        �� u�P���� u�W�        =�s� V        @�s� ub�        @�G� Pi�p� P        ���� ub����� R���� ub�        ���� P        ��² P        8�L� SL�P� �         ���� V���� ut����� tp����� V��ϳ ut�        ���� us����� to���ϳ us�        ���� R��ɳ R        ���� us���ɳ Pɳϳ us�        ��ɳ R        ��ϳ 	��        ��ɳ r�        ��ɳ Qɳϳ v�        ׳߳ Q� � Q        ��� us��� � P �� us�        � � Q        � � q�        V�#� 0�+�E� 0�E�n� 2�n��� 0�͵c� 0�        V� � 	��+��� 	��͵c� 	��        b�� V+�9� Vn��� V͵� V.�9� V        ���� P˴�� P+�H� P        ���� uS˴մ uS���� 1�        n�q� P        ��� V        {��� V͵� V.�9� V        {��� 	��͵� 	��.�9� 	��        ٵ� P.�1� P        }��� 1�        ͵� V.�9� V        ���� V        ���� P        ���� V        ��մ V        ´մ V        ȴ˴ P˴մ v        � � 1�N�c� 1�        � � VN�c� V        � � v�N�c� v�        �� v        S�n� 2�        S�_� R        S�Z� r        �.� 1�9�N� 1�        �.� V9�N� V        �.� v�9�N� v�        �#� v        ���� S���� �         ض� S�� �         ��ŷ Sܷ� S        ���� Q��ŷ �ܷ� Q        ��� �ŷܷ �        ��� �ŷܷ �        ��� Uŷܷ U        ��� �ŷܷ �        �$� S$��� � ŷܷ �         �� P�w� Ww�z� w�z��� Wŷܷ W        7�Q� UQ�Y� u p "�Y�k� P        l�t� Pŷڷ P        7�t� v|�ŷܷ v|�        H�O� PO�Q� v 8&�Q�Y� P        H�t� Sŷܷ S        H�t� Uŷܷ U        L�Q� u         L�O� PO�Q� v 8&�        Q�Y� P        Q�t� Uŷܷ U        7�l� � ���� � u��� �         7�d� �d�l� ����� �u��� �         �0� U]��� U���� ����� U�-� U-�.� �.�_� U         �4� �]�l� �u��� �         �0� �]��� ��_� �         �0� �]��� ��_� �         �0� �]��� ��_� �         �0� �]��� ��_� �         �0� �]��� ��_� �         �$� P$�0� � ]��� � �_� �         I�r� 0�r�v� Pv�0� ������ ��̼�� ���u� ����_� ��        r�}� 1�}�0� ������ ��̼� ���u� ����_� ��        r�}� 0�}�и ��ظ� ���� 1��0� ������ ��̼ڼ ���u� ����_� ��        r�}� 0�}��� ����ƺ 1�ƺ� ���#� 0�#�p� ��p��� ����0� ������ ��̼�� ���u� ����_� ��        '�0� � d��� � �_� �         '�0� �d��� ��_� �        ���� P��ո ��ظ0� ������ ��̼�� ���u� ����_� ��        �2� �2�w� Pߺ � P        �&� �&�*� QX�w� Q        ���� P��Ǹ ������ P��� ��'�8� ��ƺغ ��#�2� ��J�\� ��\��� P���� ������ P���� ���� P�.� ��        ��� Q'�:� Q:�S� ��S�d� 1�d��� Qƺߺ Q �� Q#�2� Q7�J� 1���ֻ ��ֻ0� QF�^� 6�^�u� Q��ٽ ��� � Q �1� ��1�H� Q        Źڹ Vڹ� 1�'�:� V:��� R���� 1�ƺߺ V�#� Q#�2� V2�7� R��̻ Rֻ� R�0� 1�F�^� R^�u� 6���Խ RԽ� V� � R!�1� P1�H� 1�        ��ֻ ��0� �F�^� ���� �H�_� �        ��ֻ ��0� �F�^� ���� �H�_� �        ��» P»ֻ �L�0� �LF�^� �L��Խ PH�_� �L        ��̻ Q̻ֻ ��0� �F�V� QV�^� ����� Q��� �H�_� �        ��ֻ ��0� �F�^� ���� �H�_� �        ��̻ Q̻ֻ ��0� �F�V� QV�^� �H�_� �        ��» P»ֻ �L�0� �LF�^� �LH�_� �L        ��� �        ��� �        ��Խ P        ��� �        ��� �        �0� �^�u� ��H� �        �0� �^�u� ��H� �        ��� S��0� u ^�u� u �H� S        �0� �^�j� Vj�u� ��&� V&�1� �1�=� V=�H� �        �0� �^�u� ��H� �        ��0� �^�j� Vj�u� �        ���� S��0� u ^�u� u         ��1� �        ��1� �        ��1� S        ��1� �        ��1� �        �� P��� ��ߺ � ��        ��ظ �L��_� �L�_��� V��0� �L����� �L��u� �L���_� �L�        ��ظ w|��0� w|����� w|��,� w|�.�u� w|���_� w|�        &�(� P(�*� r 8&�*�2� P        &�*� r 1�        &�*� �        &�*� �        &�(� P(�*� r 8&�        *�2� P        ��ظ �*�0� ����� ��u� ���_� �        6�E� p @K$"v @K$"+�ߺ� p @K$"v @K$"+�        ���� W        ���� �        ��� ����� �        ��� ����� �        ��� ����� �        ��� � ���� �         ���� P��� �D��d� �Dd�t� Pt�{� �#{��� P���� �D        ���� P���� � #��L� WL�O� w�O�� W��d� W���� W���� W        ��Ӿ �Ӿ� Pt��� �        ��O� V{�� V��d� V���� V        þϾ v8&�ϾӾ P        þӾ U        þӾ �        ǾϾ �        ǾϾ v8&�        ϾӾ P        ϾӾ �         �� �T        ��O� �DX�� �D��d� �D���� �D        ��پ �P�پI� SI�O� �P�X��� �P����� S��� �P���L� SL�d� �P����� S���� �P�        ��O� V��� V��d� V���� V        �.� �\        �)� �#        �8� � 8�_� V_�a� � a�~� V        �4� P8�]� Pa�}� P        �}� R        C�J� QJ�^� S^�_� vd_�a� � La�w� Qw�y� S        �2� � 8�Q� v a�}� v         �8� � 8�_� V_�a� � a�~� V        Z�_� V_�a� �         ���� P���� P        ���� R���� rP����� R        ���� Q���� q����� Q���� q����� Q���� r1����� Q        ���� r0���� r0���� r0���� r0���� r0        �� P        !�'� P'�B� �B�U� PU�Y� �        d��� T���� �`����� T���� �`�        ��� S�� �         7�K� PK��� �        ���� W���� � ���� W���� � ��� W�	� �        ���� S���� ����� S���� ���� S�	� �         ��� U�
� �        ��� V�	� �        ��� S�	� �         ��� W�	� �        &�G� �q��� ����� �        &�G� �q��� ����� �        &�G� �q��� ����� �        &�G� �q��� ����� �        &�G� Vq��� V���� ����� V        &�G� �q��� ����� �        &�G� �q��� ����� �        &�*� P*�G� � q��� � ���� �         -�G� � x��� � ���� �         -�G� �x��� ����� �        W�|� � ���� �         W�x� �x�|� ����� ����� �        ���� S�� � �         X�]� P        x�}� P        ���� �         ���� �         ���� P���� � ���� P���� � ���� P��	� �         ���� 1�        ���� P���� �         ��� P        0�<� � <�]� S]�_� � #`�_��� S        I�K� PK�_� R_�p� P���� 0����� R        l�r� Rr��� P���� P        l�r� 0�r�y� Qy�{� q�{��� Q���� Q        ���� � ���� Q���� � ���� q� �        ���� � ���� Q���� � ���� q� �        ���� � �G9%����� Q        �� P�� R�*� P8�=� 0�[�]� R        &�*� R*�<� P=�E� P        &�*� 0�*�1� Q1�3� q�3�<� Q=�]� Q        `��� � ���� P        d��� � ���� P        r��� � @F�%P�%� �        ���� � ���� S���� � 1� 0.( ���� S        ���� 0����� P��� 0�        ���� P���� P        ��� P        H�\� S\�`� �         ���� S���� �         	�� P�<� s         3�I� P        	�� px�3� Q        	��� S���� � ���� S���� � ���� S        3�Y� UY��� �L�        Y��� U���� U���� U        g�m� r �P�m�p� Qp�x� r �P�x��� �T�P����� �T�P����� �T�P�        u�x� Rx��� �T���� �T���� �T        ���� S���� � ���� S        ���� P���� �L���� P        ���� V���� ����� V        ���� W���� ����� W        ���� V        ���� P���� �L        ���� P        ��� P        �2� P        J�b� P        z��� P        ���� S���� �         �U� U���� U��� U        �:� R:�K� �K�U� R���� R���� R��� �\        ���� P���� �L        ���� V���� �        ?�`� V`�c� �        ?�a� Wa�c� �        ?�_� S_�c� �        ?�c� R        ?�b� U        v��� U���� �         v��� W���� �        ���� W�� � �        ���� V�� � �        ���� S�� � �        ���� U        1�>� PF�Y� P        <�>� P        M�f� 0�f�s� Ps��� V��� Vo��� V        ��� P        �� P�A� S_�a� S        ���� P        ���� P���� P���� P        ���� P���� p� �        ��� S�� �         ����  R����  R�        5���  Q�����  Q���  Q�        9��� �Q����� �Q�        ����  P�        ���� 0�        	���  S����  S�        	��� S���� u���� t���� S���� u���� S���� u���� S��� u�� S�� u        *��� �R���� �R�        *��� S���� u���� t���� S���� u���� S���� u���� S��� u�� S�� u        ���� 1���� 1�        ���� �R���� �R�        <��� 2���� 2�        <���  R����  R�        ���� �R����� �R��� �R�        ���� S���� u���� t���� S���� u���� S���� u�� S�� u        ���� 1����� 1��� 1�        ���� �R����� �R��� �R�        ���� �R����� �R��� �R�        ���� S���� u���� t���� S���� u���� S���� u�� S�� u        ��� 1����� 1��� 1�        ��� �R����� �R��� �R�        #��� �R����� �R��� �R�        #��� S���� u���� t���� S���� u���� S���� u�� S�� u        6��� 1����� 1��� 1�        6��� �R����� �R��� �R�        W��� �R����� �R��� �R�        W��� S���� u���� t���� S���� u�� S�� u        j��� 2����� 2��� 2�        j���  Q�����  Q���  Q�        5��� 1����� 1��� 1�        5��� �R����� �R��� �R�        [��� �R����� �R�        [��� S���� u���� t���� S���� u        n��� 2����� 2�        n��� �Q����� �Q�        9��� 1����� 1�        9��� �R����� �R�        _��� �R�        _��� S���� u���� t        r��� 1�        r��� �R�        ���� �R�        ���� S���� u���� t        ���� 1�        ���� �R�        ���� �R�        ���� S���� u���� t        ���� 2�        ����  P�        ���� �R�        ���� S���� u���� t        ���� 1�        ���� �R�        ���� �R�        ���� S���� u���� t        ���� 1�        ���� xR�        ��� xR�        ��� S���� u���� t        4��� hR�        4��� S���� u���� t        ���� P        ���� 1�         �� P         �� 1�        ���� W��-� W:�q� W        ���� R        ���� 1���-� 1�:�q� 1�        ���� 8	���-� 8	�:�q� 8	�        ���� V���� ud����� t`���� V�-� ud�:�?� V?�q� ud�        ���� V�� ud�        ���� uc��� uc�        ���� R�'� R        �� uc��'� P'�-� uc�        �'� R        �-� 	��        �'� r�        �'� Q'�-� v�        B�J� QS�k� Q        S�e� uc�e�k� Pk�q� uc�        S�k� Q        S�k� q�        ���� s����� � #����� s�        ���� �o����� P���� �o�        ���� R���� R        ���� �o����� P���� �o�        ���� R        ���� r�        ���� Q���� v�        `��� � �� � R        `��� ��� � r        `��� �        `��� �        k��� �        k��� � �� � R         �I� � I��� R         �I� �I��� r         �I� �         �I� �        �I� �        �I� � I��� R        ���� ����� S���� s����� S        0�9� �9�Y� SY�b� s�b�o� S        ���� P        ���� �         ���� ����� P        ���� ����� R        ���� � ���� pt�        ���� � #����� P        � � S �$� �         �� s��� P� � s� �$� � #�        r��� W���� u���� t���� W        o��� v����� u#����� t#����� v�        o��� S���� u���� t���� S        ���� W���� u���� t���� W        ���� v����� u#����� t#����� v�        ���� s����� u#����� t#����� s�        ��� s���� V���� u#����� t#����� V        E��� W���� u���� t���� W���� u        E��� S���� u���� t���� S        d��� W���� u���� t        d��� s����� u#����� t#�        �g� v�g�h� u#�h�i� t#�i��� v�        �f� Sf�h� uh�i� ti��� S        0�g� v�g�h� u#�h�i� t#�i��� v�        0�f� s�f�h� u#�h�i� t#�i��� s�        ���� s���$� V$�&� u#�&�'� t#�'�A� V        ��#� S#�&� u&�'� t'�A� S        ��#� s�#�&� u#�&�'� t#�        ���� 0����� P        ���� P        ���� � ���� px�        ���� � #����� P        �-� S-�1� �         �$� P$�-� s�-�1� � #�        P�|� �         P�u� �        ���� s���� V�� u#��� t#�� � V        ����
 v v <"����� v p "��� v p "�        ���� S��� S        ��� :�        ���� S��� S        ��� :�        ��� S         �L� �          �E� �        l�o� s�o��� V���� u#����� t#����� V        
�G� 0�G�J� q 4!�J�_� Q`�X� 0�X�g� 2�g��� 0�        p��� 	������ 	��        s��� V���� V        ���� P���� P��� Py��� P���� P���� P        ���� P���� P���� P        ��� P���� v        ���� V        ���� P        ���� R���� t ��B� t B�N� �PN�y� t y��� �P���� t ���� �P���� t ���� �P��� t �#� �P#�C� t C�L� �PL�s� t s�|� �P|��� t ���� R���� t ���� R���� t         ���� P��	� P	�3� �T        ����  ���X�  �g���  �����  �        ���� t ��	� R	�B� t B�N� �PN�y� t y��� �P���� t ���� �P���� t ���� �P��� t �#� �P#�C� t C�L� �PL�X� t g�s� t s�|� �P|��� t ���� t         	�3� S        �J� QJ�[� �\[��� Q���� �\���� Q���� �\���� Q���� �\��� Q�3� �\        �J� PJ�[� u �\��$�[��� P���� u �\��$����� P���� u �\��$����� P���� u �\��$���� P�	�	 u q �$�	�� P�3� u �\��$�        W�[� P���� P���� P���� P�	� P,�3� P        ���� V3�X� Vg��� V���� V        ���� 	��3�X� 	��g��� 	������ 	��        I�Q� P���� P        ���� 1�        3�Q� V���� V        ���� Vg��� V        ���� P        g��� V        y��� P        ���� �P�  ��X� �P�  g��� �P�  ���� �P�          G�J� q 4!�J�_� Q        G�_� P        G�P� R        �9� P        �9� P���� P        �%� ud�%�)� W)�*� t *�+� t+�-� t-�/� t/�2� t2�5� t5�6� t6�7� t7�9� t 9�[� ud�i��� ud����� ud�        �)� u`�)�[� Wi��� W���� W        �9� R        G�[� 4�        G�[� W        G�[� w         w��� 4�        w��� u`�        w��� u`        ���� P        ���� V        ���� v        ���� 1��� 1��+� 1�        ���� S�� S�� S        ���� s��� s��� s�        ���� s        ��� 1��� 1�+�;� 1�        ��� V�� V+�;� V        ��� v��� v�+�;� v�        ���� v        y��� P        u��� P���� P        y��� ud����� W���� t ���� t���� t���� t���� t���� t���� t���� t���� t ���� ud�        y��� u`����� W        y��� R        ���� P���� u`        ���� Q        ���� q        �� 1�B�K� 1�P�^� 1�        �� SB�D� SF�K� S        �� s�B�D� s�F�K� s�        �� s        .�B� 1�K�P� 1�^�n� 1�        .�B� VK�P� V^�n� V        .�B� v�K�P� v�^�n� v�        .�2� v        p��� 0����� 0����� 4���s� 0�        �#� 4�G�P� 4�U�c� 4�        �#� SG�I� SK�P� S        �#� s�G�I� s�K�P� s�        �� s        6�G� 4�P�U� 4�c�s� 4�        6�D� QP�T� Q        6�D� q�P�T� q�        6�:� q        ���� Q        ���� q        ���� 	����<� 	��E��� 	��        ��� 0�+�E� 0�E�S� 2�S��� 0�        ���� Q+�8� Q        ���� P<�K� P        ���� R���� q        ���� 1�        +�8� Q        ���� 1����� 1����� 1�        ���� Q���� Q        ���� q����� q�        ���� q        u��� 1����� 1�        u��� S���� S        u��� s����� s�        u�y� s        �)� S        �� s        ���� 0� �A� 0�A�O� 2�O��� 0�        	�� Q(�8� Q        �(� P<�G� P        �� R�� q        �� 1�        (�8� Q        $�(� ��          e�t� 1����� 1����� 1�        e�t� S���� S���� S        e�t� s����� s����� s�        e�i� s        ���� 1����� 1����� 1�        ���� Q���� Q        ���� q����� q�        ���� q        ���� Q        ���� q        ��� �,�i� Wl��� W���� W���� ����� W ��� W        ���� 0����� P���� p 4!����� P���� 0����� P���� 0�        �� P��� uT���� uT���� uT        ��� 	������ 	������ 	��        ��� V���� V��A� VY�b� Vg�u� V        ,�T� Pl��� P        �� �  _�b� Pb�e� vi�l� P        [�i� V���� V �� V        [�i� 	������ 	�� �� 	��        e�i� V        �<� V        i�l� P        ���� P �� P        _�e� 1�        ���� V �� V        N�i� �"�  ���� �"�   �� �"�          !�0� 1�Y�b� 1�g�u� 1�        !�0� SY�[� S]�b� S        !�0� s�Y�[� s�]�b� s�        !�%� s        C�Y� 1�b�g� 1�u��� 1�        C�Y� Vb�g� Vu��� V        C�Y� v�b�g� v�u��� v�        C�G� v        ���� 4�        ���� �Ĵ          ���� P        ���� W        ���� w        ����
 v v <"����� v p "���� v p "�        ���� S��� S        ���� :�        ���� S���� S        ���� :�        ���� S        )��� 0����� 2����� 0��� 0�        G�I� PI�g� Qg��� uT��� uT���� Q��� uT        G��� 	���� 	��        P��� S��� S���� S
�� S        _��� V���� V�Q� Vc��� V���� P        _�g� Vi��� P���� Pc�� P���� P        ?�\� ��  \�g� P���� P���� sc��� �  ���� ��          _�i� V���� P        \�g� P        ���� S        _��� �Y�  ��� �Y�  ���� �Y�          i��� Pc�� P        i��� uc�s� Qs�}� u        ���� P        ���� 1�        c�� P        c�}� u}�� Q        c��� �          ���� S�c� S        ���� 	������ V�c� 	��        ,�4� P        ���� 1�        �<� S        ���� S<�c� S        <�c� S        ���� 1����� 1�
�� 1�        ���� V���� V
�� V        ���� v����� v�
�� v�        ���� v        ���� 1���
� 1�        ���� W��
� W        ���� w���
� w�        ���� w        �� V        �
� v        )�@�
 v v <"�T�h� v p "����� v p "�        2�R� ST��� S        6��� :�        6�R� ST��� S        T��� :�        T��� S        ��� 0��-� 2�-��� 0�        ���� R��� R        �� P        ���� 1�        ��� R        �-� 2�        �'� R        �"� r        C�R� 1�y��� 1����� 1�        C�R� Sy�{� S}��� S        C�R� s�y�{� s�}��� s�        C�G� s        e�y� 1����� 1����� 1�        e�s� Q���� Q        e�s� q����� q�        e�i� q        ���� 	������ 	����	� P	�� 	���$� P$��� 	��        ���� 0���	� 0�	�$� 2�$�D� 0�W��� 0�        ���� P���� P        ��� P�#� ud#�$� t`        ���� R        ���� P        �$� 2�        �"� S        �� s        5�D� 1����� 1����� 1�        5�D� S���� S���� S        5�D� s����� s����� s�        5�9� s        m��� 1����� 1�        m�~� S���� S        m�~� s����� s�        m�q� s        ��� 0��$� 6�$��� 0�        ��#� u#�$� t$��� u        ��#� u#�$� t$��� u        ���� P        �$� 6�        �� R        �� r        :�I� 1�p�y� 1�~��� 1�        :�I� Sp�r� St�y� S        :�I� s�p�r� s�t�y� s�        :�>� s        \�p� 1�y�~� 1����� 1�        \�j� Qy�}� Q        \�j� q�y�}� q�        \�`� q        ��� 0��@� 0�@�_� 2�_��� 0�        ���� P�� P,�B� P        ���� R�(� R        ���� P�"� P"�&� rr�        �(� R        ���� u���� t ���� t        ���� R        J�_� 2�        J�V� R        J�Q� r        u��� 1����� 1����� 1�        u��� S���� S���� S        u��� s����� s����� s�        u�y� s        ���� 1����� 1����� 1�        ���� Q���� Q        ���� q����� q�        ���� q        ��� r        !�\� 0�|��� 0�        !�s� 	��|��� 	��        +�L� P|��� P        /�H� VH�L� QL�\� V|��� Q���� V        /�L� P|��� P        P�W� P        2�@� p@K$"r @K$"-�@�I� p@K$"p@K$"-�|��� p@K$"r @K$"-����� p@K$"p@K$"-����� p@K$"r@K$"-�        |��� 	��        >�H� VH�L� QL�\� V���� V        >�L� P        >�\� �4�  ���� �4�          \�s� 1�        \�o� R        \�j� r        ���� 1����� 1����� 1�        ���� S���� S���� S        ���� s����� s����� s�        ���� s        ���� 1����� 1����� 1�        ���� Q���� Q        ���� q����� q�        ���� q        �� r        =�Y� 0�`�z� 0���� 0�        =�Y� 	��`�� 	��        G�Y� P`�j� P        K�Y� P`�j� P        n�u� P        S�Y� 	��        `�j� P        z��� 1�        z��� R        z��� r        ���� 1����� 1���� 1�        ���� S���� S���� S        ���� s����� s����� s�        ���� s        ���� 1����� 1��� 1�        ���� Q���� Q        ���� q����� q�        ���� q         �u� 	��u�z� Pz�� 	��        ?�d� 0�u�z� 0�z��� 1���� 0�        H�T� P        L�T� P        ���� 1�        ���� S        ���� s        ���� 1����� 1���� 1�        ���� S���� S���� S        ���� s����� s����� s�        ���� s        ���� 1����� 1��� 1�        ���� S���� S�� S        ���� s����� s��� s�        ���� s        .�c� Sc�e� ue�h� th��� S���� u���� t���� S���� u�� � S �� u�� S�� u        s��� P        ���� 1����� 1� �� 1�        ���� V���� V �� V        ���� v����� v� �� v�        ���� v        ���� 1��� � 1��� 1�        ���� V�� � V�� V        ���� v��� � v��� v�        ���� v        3�:� r        X�e� 0�o��� 0����� 4���9� 0�        s��� P���� t ���� t        ���� 4�        ���� R        ���� r        ���� 1��� 1��)� 1�        ���� S�� S�� S        ���� s��� s��� s�        ���� s        ��� 1��� 1�)�9� 1�        ��� Q�� Q        ��� q��� q�        ���� q        Y�`� r        ~��� 0����� 0����� 4���Y� 0�        ���� P        ���� 4�        ���� R        ���� r        ��� 1�-�6� 1�;�I� 1�        ��� S-�/� S1�6� S        ��� s�-�/� s�1�6� s�        ���� s        �-� 1�6�;� 1�I�Y� 1�        �-� W6�;� WI�Y� W        �-� w�6�;� w�I�Y� w�        �� w        ���� P���� uT� �  uT        ���  	��        ���� V���� R���� uT���� tP��D  uTm �  uT� �  V� �  uT        ���� P(�/� P| �  P� �  P        s�t� uu<"�        ���� P        � �  V        � �  P        ���� P(�4� P4�0  uP        ��D   �m �   �� �   �        ���� V��D  Vm �  V� �  V        4�0  S        C�x� Qx��� uL���� Q���� uL���� Q���� uL���� Q��   uL    Q 0  uL        L�x� Px��� w uL��$����� P���� w uL��$����� P���� w uL��$����� P��   w uL��$�    P 	 	 w q �$�	   P 0  w uL��$�        ���� P���� P���� P��   P 	  P) 0  P        ��,� uT0 3  R3 D  uTm �  uT� �  uT        ��,� 	��0 D  	��m �  	��� �  	��        < D  P� �  P        �� 1�        0 D  uT� �  uT        �,� uTm �  uT        "�(� P        m �  uT        | �  P        ��D  ���  m �  ���  � �  ���          R m  2�        R ^  R        R Y  r        � A 0�A] 6�]� 0�        	 Q&8 Q        ! P<C P         R q         1�        &8 Q        & ��          K] 6�        KW R        KR r        s� 1��� 1��� 1�        s� S�� S�� S        s� s��� s��� s�        sw s        �� 1��� 1��� 1�        �� Q�� Q        �� q��� q�        �� q         B � B] S]o � o� S         9 �9> PBb �bk Po� �        .@ VBm Vo� V        4< v� fi v�         Bm Vo� V        Sn Wo� W        W�  �        Wn Wo� W        o�  �        o� W        �� ��� Q        �� r        �� R�� �        �� q        �� r  ��� R        � � ' P        �� �� R' R        
 J�        
 S � � <"�        
 s        
 	��        
 s� � � <"#�        
 Q        
 s	�� R s	��        08 �8B Q        4A � � <"�AB � r "�        4A � � <"#        PX �Xb Q        Ta � � <"�ab � r "�        Ta � � <"#        �� R        �� R R        �� u        �� ud��� Q�� t �� t�� t�� t�� t�� t�� t�� t�� ud�        �� P�� t �� t�� t�� t�� t�� t�� t        �� V�W��� V�W�L V�W�bk V�W�p~ V�W�        �� P�� ud        � W        �� w        ,; 1�bk 1�p~ 1�        ,; Sbd Sfk S        ,; s�bd s�fk s�        ,0 s        Nb 1�kp 1�~� 1�        Nb Wkp W~� W        Nb w�kp w�~� w�        NR w        � R        � RAE R        � u        �� ud��� Q�� t �� t�� t�� t�� t�  t  t t ud�        �� P�� t �� t�� t�� t�  t  t t        � V�W�( V�W�F| V�W��� V�W��� V�W�        *- P-. ud        *? W        *. w        \k 1��� 1��� 1�        \k S�� S�� S        \k s��� s��� s�        \` s        ~� 1��� 1��� 1�        ~� W�� W�� W        ~� w��� w��� w�        ~� w        3 R        3 Rqu R        7 u        ! ud�!% Q%& t &+ t+- t-. t./ t/0 t01 t13 t37 ud�        ) P)+ t +- t-. t./ t/0 t01 t13 t        .E V�W�HX V�W�v� V�W��� V�W��� V�W�        Z] P]^ ud        Zo W        Z^ w        �� 1��� 1��� 1�        �� S�� S�� S        �� s��� s��� s�        �� s        �� 1��� 1��� 1�        �� W�� W�� W        �� w��� w��� w�        �� w        ;c R        5c R�� R        ;g u        ;Q ud�QU QUV t V[ t[] t]^ t^_ t_` t`a tac tcg ud�        ;Y PY[ t [] t]^ t^_ t_` t`a tac t        ^u V�W�x� V�W��� V�W��� V�W�  V�W�        �� P�� ud        �� W        �� w        �� 1��� 1�  1�        �� S�� S�� S        �� s��� s��� s�        �� s        �� 1��  1� 1�        �� W�  W W        �� w��  w� w�        �� w        k� R        e� R�� R        k� u        k� ud��� Q�� t �� t�� t�� t�� t�� t�� t�� t�� ud�        k� P�� t �� t�� t�� t�� t�� t�� t        �� V�W��� V�W��	 V�W�"	+	 V�W�0	>	 V�W�        �� P�� ud        �� W        �� w        �� 1�"	+	 1�0	>	 1�        �� S"	$	 S&	+	 S        �� s�"	$	 s�&	+	 s�        �� s        	"	 1�+	0	 1�>	N	 1�        	"	 W+	0	 W>	N	 W        	"	 w�+	0	 w�>	N	 w�        		 w        �	�	 R        �	�	 R

 R        �	�	 u        �	�	 ud��	�	 Q�	�	 t �	�	 t�	�	 t�	�	 t�	�	 t�	�	 t�	�	 t�	�	 t�	�	 ud�        �	�	 P�	�	 t �	�	 t�	�	 t�	�	 t�	�	 t�	�	 t�	�	 t        �	�	 V�W��	�	 V�W�
<
 V�W�R
[
 V�W�`
n
 V�W�        �	�	 P�	�	 ud        �	�	 W        �	�	 w        
+
 1�R
[
 1�`
n
 1�        
+
 SR
T
 SV
[
 S        
+
 s�R
T
 s�V
[
 s�        
 
 s        >
R
 1�[
`
 1�n
~
 1�        >
R
 W[
`
 Wn
~
 W        >
R
 w�[
`
 w�n
~
 w�        >
B
 w        �
�
 R        �
�
 R15 R        �
�
 u        �
�
 ud��
�
 Q�
�
 t �
�
 t�
�
 t�
�
 t�
�
 t�
�
 t�
�
 t�
�
 t�
�
 ud�        �
�
 P�
�
 t �
�
 t�
�
 t�
�
 t�
�
 t�
�
 t�
�
 t        �
 V�W� V�W�6l V�W��� V�W��� V�W�         P ud        / W         w        L[ 1��� 1��� 1�        L[ S�� S�� S        L[ s��� s��� s�        LP s        n� 1��� 1��� 1�        n� W�� W�� W        n� w��� w��� w�        nr w        �# R        �# Rae R        �' u        � ud� Q t  t t t t  t ! t!# t#' ud�        � P t  t t t  t ! t!# t        5 V�W�8H V�W�f� V�W��� V�W��� V�W�        JM PMN ud        J_ W        JN w        |� 1��� 1��� 1�        |� S�� S�� S        |� s��� s��� s�        |� s        �� 1��� 1��� 1�        �� W�� W�� W        �� w��� w��� w�        �� w        +S R        %S R�� R        +W u        +A ud�AE QEF t FK tKM tMN tNO tOP tPQ tQS tSW ud�        +I PIK t KM tMN tNO tOP tPQ tQS t        Ne V�W�hx V�W��� V�W��� V�W��� V�W�        z} P}~ ud        z� W        z~ w        �� 1��� 1��� 1�        �� S�� S�� S        �� s��� s��� s�        �� s        �� 1��� 1�� 1�        �� W�� W� W        �� w��� w�� w�        �� w        [� R        U� R�� R        [� u        [q ud�qu Quv t v{ t{} t}~ t~ t� t�� t�� t�� ud�        [y Py{ t {} t}~ t~ t� t�� t�� t        ~� V�W��� V�W��� V�W� V�W� . V�W�        �� P�� ud        �� W        �� w        �� 1� 1� . 1�        �� S S S        �� s� s� s�        �� s        � 1�  1�.> 1�        � W  W.> W        � w�  w�.> w�        � w        �� R        �� R�� R        �� u        �� ud��� Q�� t �� t�� t�� t�� t�� t�� t�� t�� ud�        �� P�� t �� t�� t�� t�� t�� t�� t        �� V�W��� V�W��, V�W�BK V�W�P^ V�W�        �� P�� ud        �� W        �� w         1�BK 1�P^ 1�         SBD SFK S         s�BD s�FK s�         s        .B 1�KP 1�^n 1�        .B WKP W^n W        .B w�KP w�^n w�        .2 w        * P*^ V^c �P�        * R*] S        * Q*c �\        * Q*2 w p �2a W        *6 PAN P        �� 0��� S�� � �� 0�        �� P�� P        �� � �� S�� �         � 0�"} 0�        �! u!" �"e uef tf} u        Ef 0�        �� 0��� P�� 0��� S�� P        5� 0��� S�� � �� 0�        5m � m� S�� � �� S�� �         ?Z 0�Ze Pv} P}� 0�        �� P� P        @O 0�Os Ssu Pu� 0��� P         
 �         ,A P        �� s��� � #��� s�        �� �o��� P�� �o�        �� R�� R        �� �o��� P�� �o�        �� R        �� r�        �� Q�� v�         S  �         H\ S\` �         �� S�� �         �� S�� �         ": s�:< � #�<` s�        %T �o�TZ PZ` �o�        %- R<Z R        <T �o�TZ PZ` �o�        <Z R        <Z r�        CZ QZ` v�        x� S�� �         �� S�� �         � S �         �� P�\ W^� W        �� S        �� P�[ V^� V        �� 0�        �� P�| W~� W        � S�� S        �� P�{ V~� V         P� W� W        � S� S        )3 P3� ud�� t`�� ud        SV PV� p��� p��� p��� p�        / �        �� P�� V        �� S        �� ud        �� S        �!�! S�!�! �         �!�! ��~        ["x" Sx"{" t	��{"" t	��"�" t	���"�" t	���"�" t	���"�" S        t"~" P~"�" V�"�" P        �"�" ��"�" �#;# �#�;#C# ��#�# U        �"�" � �"�" s��"]# Sa#�# S        �"# V#^# Va#�# V        �"_# W_#a#
 � �"1�a#�# W        #G# R        �#�# P        �#�# S�# $ �         ($<$ S<$@$ �         \$b$ p�b$�$ u#��$% u#�(%�% u#��%�% u#�        s$�$ P�$�$ u#�$�$ P�$�$ u#(%3% P3%B% u#E%S% PS%b% u#h%s% Ps%�% u#        s$�$ Q�$�$ Q(%B% QE%b% Qh%�% Q        s$�$ ud��$�$ P�$�$ ud�(%�% ud�        }$�$ ud�$�$ p �$�$ ud(%B% udE%b% udh%�% ud        �$�$ �	�        �$�$ ud��$�$ P�$�$ ud�        �$�$ �	�        �$�$ ud��$�$ P�$�$ ud�        (%E% % 	�        (%3% ud�3%B% PB%E% ud�        E%h%  	�        E%S% ud�S%b% Pb%h% ud�        h%�% �	�        h%s% ud�s%�% P�%�% ud�        �%�% Q�%�% Q        �%�% uc��%�% R�%�% uc�        �%�% Q        �%�% q�        �$�$ ud�%% S        �$�$ uc�%% uc�        �$�$ R%% R        �$�$ uc��$�$ Q�$�$ uc�        �$�$ R        �$�$ 	��        �$�$ r�        �$�$ Q�$�$ s�        �%& u&	& t	&,& u,&/& t/&Q& uQ&T& tT&|& u|&& t&�& u�&�& t�&�& u�&�& u        �%�% s 	&& s /&?& s T&j& s &�& s         �%	& �	�        �%& u&	& t        T&& % 	�        T&|& u|&& t        	&/&  	�        	&,& u,&/& t        5&T& �	�        5&Q& uQ&T& t        &�& �	�        &�& u�&�& t        �&�& u�&�& u        �&�& Q�&�& Q        �&�& ug��&�& R�&�& ug�        �&�& Q        �&�& q�        h(|( S|(�( �         �(�( S�(�( ��(�( S�(�( �        N)Z) Q        N)Z) R        N)Z) P        �)�) � �)�) [        �)�) S�)�) �             $    P$   R    VR   U    �P�U   h    Ph   t    Vt   �    P�   �    �P�        $   P    V        >   P    W        �   �    P�   �    �P�        �   �    V�   �    P        �   �    Q        �   �    R           	   P	     S     �P�  @   S@  B   �P�B  [   S              R  9   P9  =   Q=  B   �R�B  [   P        	     R  9   P9  =   Q=  >   �R�>  [   P          -   RB  Y   R        $  -    �-  =   RB  [   O�        `  j   Pj  k   �P�k  �   P�  �   �P��  c   Pc  n   �P�n     P  
   �P�
  +   P        `  �   R�  �   �R��  �   R�  n   �R�n  t   Rt     �R�  +   R        �  �   S�     S  B   SF  j   Sn  �   S
     S  +   S        �  �   q ���  �   p3%1��  �   Qt  �   Q
     Q        �  �    -	��  �   Rt  �   R
     R        �  �   �-	�t     �-	�        �  �   p        �  
   Q     Q        �  
   V     V        �  
   V        �  
   Q        �     P  
   �P�        �  
   R        �  �   W�  �   �h        �  �   V�  �   r�  �   V�  �   �d        �  �   P        �  �   W        �  �   0��     R  &   Q&  <   R<  n   Qn  t   0�          &   Q&  +   R:  S   Q        0  =   P=  Y   VY  [   �P�[  �   V        0  =   R=  Z   WZ  [   �R�[  �   W        0  =   Q=  �   �Q�        �  �   P�  �   �P��  �   P�     �h        �  �   R�  �   �R��  �   R�     �R�        �  �   P�     �h          $   0�a  �   1�          s   Rs  ~   p �  �   R        $  4   0�4  W   SW  Y  	 s u 'w "�\  a   P        �  �   P�  �   pt��  �   �P��  �   P�  �   �P��  �   P�  �   �P�        �  �   S�  �   P�  �   S�  �   rr1$"2$q "�        �  �   P�     S     �P�  )   S)  *   �P�*  /   S        	     p�"  *   P*  -   p�-  /   P        0  :   P:  ;   �P�;  N   PN  ~   S~  �   �P��  �   S�  �   �P�        O  }   P}  �   r�  �   P        W  }   P}  �   r        W  ~   S~  �   �P�        n  �   R        �  �   P�  �   �P��  �   P�  �   pt��  �   �P�        �  �   P�  �   p  �        �  �   P�     S  !   �P�!  �   S        �  �   P�     V!  z   Vz  �   P�  �   V        �  �   P�     V!  z   V�  �   V        �     S!  z   S�  �   S        �     W!  z   W�  �   W        @  z   w�        �  �   P�  �   S�  �   �P��     S        �  �   R�  �   R�  �   �R��  �   R�     R           -   P-  �   �P��  �   P�  �   �P�        2  �   R        2  B   PB  e   q#e  g   Pg  �   q#        2  \   P_  r   Ps  �   P        �  �   P�  �   �P�        �  �   P�  �   V�  �   �P��  	   V	  		   �P�        �  �   R�  		   �R�        �  �   P�  		   P        	  g	   �g	  �	   W�	  �	   �        	  g	   �g	  �	   V�	  �	   �        	  0	   �0	  2	   V2	  4	   �4	  e	   Ve	  g	   �g	  �	   V        	  4	   �4	  f	   Wf	  g	   �g	  �	   W        %	  )	   Pg	  �	   P�	  �	   P        g	  �	   P�	  �	   P        {	  �	   2��	  �	   S�	  �	   2�        �	  �	   P�	  �	   P        �	   
   P 
  �
   V�
  �
   �P�        �	   
   R 
  
   S
  �
   �R�        
  
   P        
  
   S
  �
   �R�        
  �
   V�
  �
   �P�        
  
   0�
  %
   s �R�;
  ~
   s �R�        
  %
   RD
  g
   Rg
  ~
   �_        
  ;
   VD
  ~
   V        J
  ~
   V        �
  �
   P�
  D   SD  H   �P�        �
  �
   R�
  H   �R�        �
  G   UG  H   �G�        �
  D   SD  H   �P�        �
  �
   P        �
  G   UG  H   �G�        �
  D   SD  H   �P�        �
  �
   0��
  8   V        �
  �
   Q�
     Q  8   ��        �
  �
   S�
  8   S           8   S        P  o   Po  T   ST  X   �P�X  �   S�  �   �P��  �2   S        P  �   R�  L   u�L  X   �R�X  [   R[  �   u��  �   t��  �   R�  -   u�-  :   R:  h   u�h  p   Rp  d   u�d  k   Rk  �   u��  �   R�  �   u��  �   R�  3   u�3  C   RC  �   u��  �   R�  3   u�3  C   RC  �   u��  �   R�     u�  �   �R��  �   R�     u�  	   R	  1   u�1  >   R>  T   u�T  }   R}  �   u��  �   �R��  �   R�  �   u��  �   R�  #   u�#  >   R>  �   �R��  �   R�  #   u�#  0   R0  �   u��  �   R�     u�  "   R"  f   u�f  �   R�  �   u��     R  �   u��     R  �   u��  �   R�  �   u��     R  7   u�7  U   RU  y   u�y     R  �   u��  �   R�  �   u��  �   R�  �   u��  �   R�  �   u��  �   R�     u�     R  3   u�3  :   R:  n   u�n  u   Ru  �   u��  �   R�  �   u��  �   R�  �   u��  �   R�  �   u��     R  s   u�s  v   Rv  �   u��  �   R�  Y   u�Y  t   Rt  �   u��  �   R�  S   u�S  ^   R^  �   u��  �   R�     u�  G   RG  �   u��  �   R�  /   u�/  @   R@  �   u��  �   R�  �   u��  �   R�      u�       R   /    u�/   6    R6   P    u�P   m    Rm   �    u��   �    R�   !   u�!  !   R!  4!   u�4!  C!   RC!  �!   u��!  _"   �R�_"  &$   u�&$  -$   R-$  �$   u��$  s%   �R�s%  �%   u��%  &   R&  }&   u�}&  �&   R�&  �&   u��&  �&   �R��&  �&   R�&  g'   u�g'  �'   R�'  (   u�(  '(   �R�'(  J(   RJ(  )   u�)  1)   R1)  f)   u�f)  )   �R�)  *   u�*  !*   R!*  �*   �R��*  ,   u�,  ,   R,  X-   u�X-  t-   �R�t-  F.   u�F.  x.   �R�x.  p/   u�p/  �/   R�/  F0   u�F0  q0   �R�q0  �0   u��0  �0   �R��0  �0   R�0  /1   u�/1  D1   RD1  S1   u�S1  }1   �R�}1  �1   u��1  �1   R�1  �1   �R��1  �1   u��1  2   R2  C2   u�C2  �2   �R��2  �2   u�        P  �   Q�  L   u�X  [   Q[  �   u��  �   �Q��  �   Q�  -   u�-  8   Q8  h   u�h  v   Qv  �   u��  d   u�d  o   Qo  �   u��  �   Q�  �   u��  �   Q�  3   �Q�3  C   QC  �   �Q��  �   Q�  3   �Q�3  C   QC  �   �Q��  �   Q�     u�  �   �Q��  �   Q�     �Q�     Q  1   �Q�1  <   Q<  T   u�T  z   Qz  �   �Q��  �   Q�  �   u��  �   Q�  #   �Q�#  0   Q0  >   u�>  �   �Q��  �   Q�  #   �Q�#  )   Q)  d   u�d  �   �Q��  �   Q�     u�  "   Q"  f   �Q�f  �   Q�  �   �Q��  )   Q)  �   u��     Q     u�  �   �Q��  �   Q�  �   u��     Q  M   u�M  7   �Q�7  U   QU  y   u�y  �   Q�  �   u��  �   Q�  �   u��  �   Q�  �   u��  �   Q�  �   u��  �   Q�     u�     Q  3   u�3  >   Q>  n   u�n  y   Qy  �   u��  �   Q�  �   u��  �   Q�  �   u��  �   Q�  �   u��     Q  s   �Q�s     Q  �   u��  �   Q�  Y   u�Y  t   Qt  �   �Q��  �   Q�  S   �Q�S  \   Q\  �   u��  �   �Q��  �   Q�     �Q�  E   QE  U   u�U  �   �Q��  �   Q�  /   �Q�/  @   Q@  e   �Q�e  �   u��  �   Q�  �   u��  �   Q�      u�       Q   /    u�/   :    Q:   P    u�P   m    Qm   �    u��   �    Q�   !   �Q�!  !   Q!  4!   u�4!  C!   QC!  x!   u�x!  �!   u��!  $   �Q�$  $   u�$  &$   P&$  -$   Q-$  �%   �Q��%  �%   u��%  &   Q&  }&   �Q�}&  �&   Q�&  �&   u��&  �&   �Q��&  �&   Q�&  g'   �Q�g'  o'   Qo'  '(   �Q�'(  G(   QG(  )   u�)  1)   Q1)  )   �Q�)  *   u�*  !*   Q!*  +   �Q�+  +   u�+  v+   �Q�v+  �+   Q�+  �+   �Q��+  ,   u�,  @,   Q@,  o,   u�o,  �,   �Q��,  �,   Q�,  -   u�-  #-   �Q�#-  X-   u�X-  t-   �Q�t-  �-   u��-  �-   Q�-  F.   u�F.  p/   �Q�p/  }/   Q}/  �/   u��/  0   �Q�0  F0   u�F0  q0   �Q�q0  �0   u��0  �0   �Q��0  �0   Q�0  �1   �Q��1  �1   u��1  �1   Q�1  �1   �Q��1  �1   u��1  2   �Q�2  C2   u�C2  �2   �Q��2  �2   Q�2  �2   u�        P  L   0�X  �   0��  �   Q�  $   0�$  #-   0�#-  X-   QX-  �2   0�        w  {   Q{  �   u�@  �   u�o&  }&   u�-  X-   u�        P  L   0�X  w   0�w  �   1��  @   0�@  �   V�  $   0�$  $   V$  o&   0�o&  }&   V}&  -   0�-  X-   VX-  �2   0�        �  �   0��  L   V�+  ,   V�,  �,   V�,  -   v��-  �-   V2  C2   V�2  �2   V        �  L   (��+  ,   (��-  �-   (�        �  L   S�+  ,   S�-  �-   S        �+  ,   S          L   )��+  �+   )��-  �-   )�          L   S�+  �+   S�-  �-   S        �+  �+   S        X  t   Pt  {   r|�|  �   P�  �   p�  �   P7  e   Po&  }&   P'(  �(   P�(  �(   u�~)  )   P-  )-   P�1  �1   u�~        |  �   P�  �   p�  �   P)  )   P        X  �   S8(  )   S�1  �1   S        X  t   Pt  {   r|�|  �   P�  �   p�  �   P8(  �(   P�(  �(   u�~)  )   P�1  �1   u�~        X  [   0�8(  L(   0�L(  e(   Q        �  �   R        �  �   P�  �   p�  �   P        e(  �(   P�(  �(   u�~)  )   P�1  �1   u�~        e(  )   S�1  �1   S        w(  �(   R�(  �(   r|�        �(  �(   W�(  �(   s��(  �(   Q�1  �1   Q        �(  �(   R�(  �(   V�1  �1   R        �(  �(   R�(  �(   V�1  �1   R        �  �   S�  �   �P�        �  �   0��  �   u��!  �!   P$  &$   0�        w  �   P�1  �1   P        �  �   P�  �   P$  $   P        �  d   Wx!  �!   W$  &$   W        �    	 v 6	�#  d  	 v 6	�        �     P,  L   PL  d   u�        �  #   S,  d   Sx!  �!   S        :  d   S        �  �  	 v �6	��  3  	 v �6	�        �  �   R�     R  3   u�        �  �   S�  3   S�"  #   S        	  3   S        C  U  	 v �6	�s  �  	 v �6	�        C  U   R{  �   R�  �   u�        C  s   S{  �   S�!  �!   S        �  �   S        �  �  	 v h6	��  3  	 v h6	�        �  �   R�     R  3   u�        �  �   S�  3   S�!  �!   S        	  3   S        C  U  	 v M6	�s  �  	 v M6	�        C  U   R{  �   R�  �   u�        C  s   S{  �   S�"  �"   SD+  v+   S        �  �   S        �  �   u�#�  �   t �  �   t�  �   t        �  �   S        �  �   u�        �  �   S              w q �  �   W        �  �   u��        �  �   S              0�  �   V          %   RK  k   Rk  �   u�          ?   SK  �   S        Y  �   S        �  �  	 v �5	��    	 v �5	�        �  �   R�  �   R�     u�        �  �   S�     S�#  �#   S        �     S        	     Rv+  �+   R�+  �+   u�        	  1   Sv+  �+   S        �+  �+   S        e  �   Wg'  t'   Wt'  (   u�)  )   Wo,  �,   u��0  �0   W/1  S1   u�}1  �1   u��1  2   u�        e  �   u�g'  (   u�)  f)   u�o,  �,   u��0  �0   u��0  �0   u�/1  M1   u�R1  S1   u�}1  �1   u��1  
2   u�#        e  �   0�g'  |'   0�|'  �'   V�'  �'   u�)  )   0��0  �0   0�        �'  '(   (�R1  �1   (�        �'  '(   SR1  �1   S        }1  �1   S        �'  '(   )�R1  }1   )�        �'  '(   SR1  }1   S        R1  }1   S        )  )   (��0  �0   (�        )  )   S�0  �0   S        �0  �0   S        U)  )   )��0  �0   )�        U)  )   S�0  �0   S        �0  �0   S        �  �  	 v 6	��  #  	 v 6	�        �  �   R�     R  #   u�        �  �   S�  #   S_"  q"   S        �  #   S        .  9   P9  >   Q>  �   u��!  �!   u��&  �&   u�F0  G0   u�        3  �   W�!  �!   W�&  �&   WF0  q0   W        3  �   6	��!  _"   6	��&  �&   6	�F0  q0   6	�        3  �   S�!  _"   S�&  �&   SF0  q0   S        3  �   8��!  _"   8��&  �&   8�F0  q0   8�        3  >   0�>  E  	 v 6	�c  �  	 v 6	�        >  E   Rk  �   R�  �   u�        >  c   Sk  �   S�!  _"   S�&  �&   SF0  q0   S        y  �   S        �!  �!   w p ��!  �!   W        �!  _"   S        �!  �!   0�        �!  "   R'"  G"   RG"  _"   u�        �!  "   S'"  _"   S        5"  _"   S        �&  �&    �F0  q0    �        �&  �&   SF0  q0   S        F0  q0   S        �  �  	 v 6	��  #  	 v 6	�        �  �   R�     R  #   u�        �  �   S�  #   Sq"  �"   S        �  #   S        �#  �#   V�#  $   v�        �#  $   W        W  d   0�d  u  	 w 6	��  �  	 w 6	�        d  u   P�  �   P�  �   u�        d  �   S�  �   S�#  $   S        �  �   S        )  �)   S        �  �   Q        �     V        f  u   S        �  �  	 v >6	��  �  	 v >6	�        �  �   R�  �   R�  �   u�        �  �   S�  �   S�"  �"   S        �  �   S        �     S             u�          7   RC!  `!   R`!  d!   v �-  �-   R�-  �-   v         (  3   W3  �   u��0  /1   u�        (  �   u��0  /1   u�        (  D   rD  �   u��0  �0   r�0  /1   u�        +  .   P.  D   rD  �   u��0  �0   r�0  /1   u�           O   WO     u��*  +   u�0  40   W        &  O   1�O     V�*  +   V0  40   1�        &  O   WO  �   P�*  +   P0  40   W        �*  +   S        �  s   W&$  �$   W�$  �$   t            	 v \6	�3  s  	 v \6	�             R;  [   R[  s   u�          3   S;  s   S        I  s   S        -$  5$  	 v a6	�O$  �$  	 v a6	�        -$  5$   RW$  w$   Rw$  �$   u�        -$  O$   SW$  s%   SF.  x.   S        e$  �$   S        �$  �$   W�$  �$   t        �$  s%   SF.  x.   S        �$  s%   u�F.  x.   u�        �$  s%   SF.  x.   S        �$  �$   w u���$  s%   WF.  x.   W        �$  s%   u��F.  x.   u��        �$  s%   SF.  x.   S        �$  �$   0��$  O%   V        �$  �$   R%  7%   R7%  O%   u�        �$  %   S%  O%   S        %%  O%   S        O%  s%   }�F.  x.   }�        O%  s%   SF.  x.   S        F.  x.   S        �  �   V        �  �   P�  �   Q�)  �)   P�)  *   P        �)  *   R        �)  �)   P        �)  �)   P�)  �)   P        �  �   W�  Y   u�t-  �-   u�p/  x/   Wx/  �/   u�        �  �   P�  �   s�#p/  �/   P�/  �/   s�#        �  �   P�  �   s��  Y   u�t-  �-   u�p/  �/   u�        b  r   Wr  t   u�#        b  t   V        b  �   S        b  t   0�        t  �   R�  �   R�  �   u�        t  �   S�  �   S        �  �   S        �  �  	 v �5	�  S  	 v �5	�        �  �   R  ;   R;  S   u�        �     S  S   S�#  �#   S        )  S   S        �  �   Q+  +   Q+  ?+   u�?+  D+   Q        �  �   W�  �   u�#        �  �   V        �     S        �  �   0�        �  �   R�     R     u�        �  �   S�     S        �     S        2  5   P5  �   u�x.  p/   u��/  0   u��1  �1   u�        8  �   Wx.  �.   W�.  �.   s�#�.  %/   u��/  0   W�1  �1   W        2  U   0�U  �   Vx.  p/   V�/  0   V�1  �1   V        �  �   S        �.  /   Q/  /  	 s�<#�1  �1   Q        �  �   W�  �  	 u�##        �  �   V        �  /   S        �  �   0�        �  �   R�     R  /   u�        �  �   S�  /   S          /   S        c   m    Wm   �    R�)  �)   R�1  �1   W�1  �1   s�        �   �   	 v �5	��   !  	 v �5	�        �   �    R�   �    R�   !   u�        �   �    S�   !   S#  �#   S        �   !   S        4!  C!   S        �"  �"   )�D+  v+   )�        �"  �"   SD+  v+   S        D+  v+   S        #  �#   �4	�        #  �#   S        #  �#   5�        #  !#   0�!#  5#  	 v �4	�O#  �#  	 v �4	�        !#  5#   RW#  w#   Rw#  �#   u�        !#  O#   SW#  �#   S        e#  �#   S        �%  �%  	 v 6	��%  �%  	 v 6	�        �%  �%   R�%  �%   R�%  �%   u�        �%  �%   S�%  �%   S        �%  �%   S        �%  
&   W
&  &  	 u�##        �%  &   V        �%  o&   S        �%  &   0�        &  &   R7&  W&   RW&  o&   u�        &  /&   S7&  o&   S        E&  o&   S        �&  '  	 v �5	�'  _'  	 v �5	�        �&  '   R''  G'   RG'  _'   u�        �&  '   S''  g'   S        5'  _'   S        *  !*   p        *  !*   V        *  �*   SX-  t-   S�1  �1   SC2  �2   S        *  �*   VX-  t-   V�1  �1   VC2  d2   V        *  �*   WX-  t-   W�1  �1   WC2  �2   W        !*  D*   R�*  �*   R�*  �*   u�        !*  S*   S�*  �*   S        �*  �*   S        {*  �*   0��*  �*   p r "��*  �*   R        �*  �*   P�*  �*   u��*  �*   P�*  �*   u�X-  t-   u�C2  n2   u�        �*  �*   P�*  �*   Po-  t-   P        d2  �2   S        f2  �2   S        q0  �0   Q        y0  �0   S        �2  3   P3  ,3   S,3  73   P73  83   �P�83  F3   PF3  �3   S�3  �3   P�3  E4   SE4  V4   PV4  �4   S�4  �4   P�4  E5   SE5  e5   Pe5  �5   S�5  �5   �P��5  �5   P�5  A6   SA6  _6   P_6  �6   S�6  �6   P�6  �6   S�6  �6   P�6  �6   S�6  �6   P�6  %7   S%7  67   P67  �7   S�7  �7   P�7  9   S9  /9   P/9  x9   Sx9  �9   P�9  :   S        �2  3   R3  ,3   W,3  73   R73  83   �R�83  M3   RM3  �3   W�3  �3   R�3  E4   WE4  ]4   R]4  �4   W�4  �4   R�4  E5   WE5  V5   RV5  �5   W�5  �5   �R��5  �5   R�5  A6   WA6  m6   Rm6  �6   �R��6  �6   R�6  %7   W%7  =7   R=7  �7   W�7  �7   R�7  �8   W�8  �8   R�8  �9   W�9  �9   R�9  �9   W�9  �9   R�9  :   �R�        �2  3   Q3  ,3   U,3  83   �Q�83  M3   QM3  �3   U�3  �3   Q�3  �3   U�3  �3   Q�3  E4   UE4  ]4   Q]4  �4   U�4  �4   Q�4  E5   UE5  e5   Qe5  �5   U�5  �5   �Q��5  �5   Q�5  A6   UA6  m6   Qm6  �6   U�6  �6   Q�6  %7   U%7  =7   Q=7  �7   U�7  �7   Q�7  �8   U�8  �8   Q�8  9   U9  /9   Q/9  x9   Ux9  �9   Q�9  �9   U�9  �9   Q�9  �9   U�9  �9   Q�9  :   U         3  ,3    ��8  9    �         3  3   P3  ,3   S�8  9   S        �8  9   S        M3  U3  	 v  7	�s3  �3  	 v  7	�        M3  U3   R{3  �3   R�3  �3   �_        M3  s3   S{3  �3   Se8  �8   SF9  x9   S        �3  �3   S        �3  �3  	 v �6	�4  E4  	 v �6	�        �3  �3   R4  ,4   R,4  E4   �_        �3  4   S4  E4   S        4  E4   S        ]4  e4  	 v �6	��4  �4  	 v �6	�        ]4  e4   R�4  �4   R�4  �4   �_        ]4  �4   S�4  �4   S        �4  �4   S        �4  �4  	 v �6	�5  E5  	 v �6	�        �4  �4   R5  ,5   R,5  E5   �_        �4  5   S5  E5   S        5  E5   S        E5  v5    �9  F9    �        E5  e5   Pe5  v5   S9  /9   P/9  F9   S        9  /9   P/9  F9   S        v5  �5   &��8  �8   &�        v5  �5   S�8  �8   S        �8  �8   S        �5  �5    �x9  �9    �        �5  �5   P�5  �5   Sx9  �9   P�9  �9   S        x9  �9   P�9  �9   S        �5  �5   0��5  �5  	 v �6	��5  A6  	 v �6	�        �5  �5   R6  (6   R(6  A6   �_        �5  �5   S6  A6   S        6  A6   S        Y6  �6   *��9  :   *�        Y6  _6   P_6  �6   S�9  :   S        �6  �6  	 v �6	��6  %7  	 v �6	�        �6  �6   R�6  7   R7  %7   �_        �6  �6   S�6  %7   S        �6  %7   S        =7  E7  	 v �6	�c7  �7  	 v �6	�        =7  E7   Rk7  �7   R�7  �7   �_        =7  c7   Sk7  �7   S        q7  �7   S        �7  �7    ��9  �9    �        �7  �7   P�7  �7   S�9  �9   S        �9  �9   S        �7  e8   �6	�        �7  e8   S        �7  e8   3�        �7  �7   0��7  8  	 v �6	�#8  e8  	 v �6	�        �7  8   R+8  L8   RL8  e8   �_        �7  #8   S+8  e8   S        18  e8   S        |8  �8   )�F9  x9   )�        |8  �8   SF9  x9   S        F9  x9   S        �=  �=   P�=  c>   Sc>  g>   �P�g>  b@   S        �=  �=   R�=  d>   Vd>  g>   �R�g>  �?   V�?  @   R@  b@   V        �=  �=   1�g>  k?   1��?  @   1�@  0@   0�        �=  �=   0�@  0@   0�        �=  �=   Pg>  s>   P        �>  �>  	 u U6	��>  �>  	 u U6	�        �>  �>   R�>  �>   R�>  �>   �_        �>  �>   S�>  k?   S        �>  �>   S        ?  k?   )�        ?  k?   S        <?  k?   S        �=  >    �0@  b@    �        �=  >   S0@  b@   S        >  g>   [�k?  �?   [�        >  c>   Sc>  g>   �P�k?  �?   S        �?  �?   S        @>  g>   ]�k?  �?   ]�        @>  c>   Sc>  g>   �P�k?  �?   S        k?  �?   S        p@  �@   P�@  �@   S�@  dA   �\dA  B   �P�B  iB   �\iB  dC   �P�dC  �C   �\        p@  �@   R�@  	B   W	B  B   �R�B  �C   W        �@  �@   0�_A  �A   0�B  B   0�B  )B   1�        �@  �@   0��@  -A   1�_A  �A   0�B  )B   0�dC  �C   1�        �@  �@   V�@  �@   P_A  dA   PB  B   P        rB  �B   �\2C  dC   �\        �@  -A    �dC  �C    �        �@  -A   SdC  �C   S        'A  _A   (�/B  �B   (�2C  dC   (�        'A  _A   S/B  �B   S2C  dC   S        -A  _A   S        �A  B   (��B  2C   (�        �A  B   S�B  2C   S        �B  �B   S        �A  B   )��B  2C   )�        �A  B   S�B  2C   S        �B  2C   S        rB  �B   )�2C  dC   )�        rB  �B   S2C  dC   S        2C  dC   S        �C  �C   P�C  �C   S�C  �C   �P��C  �D   S�D  �D   �P��D  �E   S        �C  �C   R�C  �C   W�C  �C   �R��C  �D   W�D  �D   �R��D  �E   W         D  �D   W�D  �D   �R��D  �E   W         D  �D   S�D  �D   �P��D  �E   S        3D  E   <�GE  wE   <��E  �E   <�        3D  �D   S�D  �D   �P��D  E   SGE  wE   S�E  �E   S        �D  �D   S        oD  �D   >��D  E   >�        oD  �D   S�D  �D   �P��D  E   S        �D  E   S        E  GE    �wE  �E    �        E  GE   SwE  �E   S        wE  �E   S        GE  wE    ��E  �E    �        GE  wE   S�E  �E   S        �E  �E   P�E  �E   �P��E  F   PF  mF   SmF  wF   �P�        �E  �E   R�E  �E   �R��E  �E   R�E  wF   �R�        �E  �E   Q�E  �E   �Q��E  F   QF  wF   �Q�        �E  �E   R�E  wF   �R�        �E  F   QF  wF   �Q�        �E  F   PF  mF   SmF  wF   �P�        �E  F   WF  F   r        �E  F   V        �E  F   PF  mF   SmF  wF   �P�        �E  F   0�        F  F   R3F  TF   RTF  mF   �o        F  +F   S3F  mF   S        9F  mF   S        �F  �F   P�F  G   UG  G   �P�G  G   UG  !G   P!G  "G   �P�"G  �G   S        �F  �F   R�F  "G   �X"G  XG   RXG  �G   �X        �F  �F   Q�F  G   �Q�G  !G   Q!G  "G   �Q�"G  XG   QXG  rG   �\rG  �G   �Q�        �F  G   0�G  "G   1�"G  �G   0�        �F  G   (�"G  �G   (�        �F  G   UG  G   �P�"G  �G   S        8G  rG   S        �F  G   )�rG  �G   )�        �F  G   UG  G   �P�rG  �G   S        �G  �G   P�G  �G   �P��G  �G   P�G  �H   V�H  �H   �P��H  �H   V�H  �H   �P��H   I   V        kH  yH   P�H  �H   P        H  H   PH  tH   W�H  �H   W�H  I   PI   I   W        H  #H   ;�#H  tH   U�H  �H   <�I   I   U        #H  [H   RI   I   R        �H  �H   0�        �H  �H   V        �H  �H   P        n  n   Pn  Dn   SDn  Hn   �P�Hn  o   So  o   �P�o  #�   S        n  #n   p #n  'n   sHn  ]n   p         *n  En   V�n  o   V�s  �s   V        `n  �n   So  �s   S�s  #�   S        `n  �n   Uo  �s   U�s  #�   U        dn  �n   Ro  $o   R$o  <o   v Hp  fp   R�p  �p   R�p  �p   v �q  �q   R�q  r   Rt  t   v ct  it   v �t  �t   R؍  �   R        �n  �n   0��n  �n   W�t  �t   0��t  �t   P        Bo  Jo   PJo  p   t p  p   �Pp  !p   t !p  Dp   �PDp  Hp   t �p  �q   t �q  �q   �P�q  �q   t r  �r   t �r  s   �Ps  js   t js  �s   �P�s  �s   t �s  �s   t �s   t   �P t  t   t Gt  ct   t �t  �t   t �t  �t   �P�t  �t   t �t  �t   �P�t  ,u   t ,u  @u   �P@u  �u   t �u  v   �Pv  �v   t �v  �v   �P�v  Rw   t Rw  fw   �Pfw  �w   t �w  �w   t �w  �w   �P�w  �x   t �x  �x   �P�x  �x   t �x  �x   �P�x  ky   t ky  }y   �P}y  �y   t �y  �y   �P�y  z   t z  #z   �P#z  az   t az  sz   �Psz  �z   t �z  {   �P{  C{   t C{  V{   �PV{  �{   t �{  |   �P|  2|   t 2|  E|   �PE|  r|   t r|  �|   �P�|  �|   t �|  �|   �P�|  \}   t \}  o}   �Po}  |}   t |}  �}   �P�}  �}   t �}  �}   �P�}  �}   t �}  �}   �P�}  �~   t �~  �~   �P�~     t   "   �P"  R   t R  a   �Pa  �   t �  
�   �P
�  �   t �  -�   �P-�  ��   t ��  ��   �P��  ƀ   t ƀ  ؀   �P؀  �   t �  &�   �P&�  /�   t /�  >�   �P>�  C�   t C�  R�   �PR�  r�   t r�  ��   �P��  �   t �  �   �P�  "�   t "�  5�   �P5�  m�   t m�  ��   �P��  ��   t ��  1�   �P1�  C�   t C�  X�   �PX�  ��   t ��  ��   �P��  �   t �  ��   �P��  �   t �  �   �P�  �   t �  0�   �P0�  P�   t P�  w�   �Pw�  ��   t ��  ��   �P��  �   t �  ��   �P��  f�   t f�  ��   �P��  ��   t ��  ��   �P��  ��   t ��  �   �P�  �   t �  #�   �P#�  (�   t (�  7�   �P7�  W�   t W�  |�   �P|�  ��   t ��  ��   �P��  Ն   t Ն  �   �P�  �   t �  �   �P�  E�   t E�  Y�   �PY�  ��   t ��  ��   �P��  �   t �  G�   �PG�  Y�   t Y�  l�   �Pl�  ��   t ��  ��   �P��  ��   t ��  ڈ   �Pڈ  '�   t '�  :�   �P:�  G�   t G�  Z�   �PZ�  _�   t _�  r�   �Pr�  ��   t ��  ��   �P��  ��   t ��  
�   �P
�  ��   t ��  ��   �P��  ��   t ��  ��   �P��  Ҋ   t Ҋ  ؊   �P؊  �   t �  ��   �P��  -�   t -�  D�   �PD�  r�   t r�  ��   �P��  ��   t ��  Ƌ   �PƋ  ��   t ��  �   �P�  ��   t ��  ��   �P��   �   t  �  �   �P�  %�   t %�  <�   �P<�  ��   t ��  ��   �P��  ؍   t �  �   t �  �   �P�  [�   t [�  a�   �Pa�  ގ   t ގ  ��   �P��  �   t �  (�   �P(�  h�   t h�  z�   �Pz�  ��   t ��  ��   �P��  ��   t ��  ��   �P��  
�   t 
�  #�   �P        6o  uo   0��p  q   0�r  *r   0�*r  1r   V7r  Rr   �TGt  Vt   �T�t  �t   0��t  �t   �T        �p  q   t #q  )q   P7r  :r   p:r  Ur   P�s  �s   PZu  ]u   P        p  -p   Q�t  �t   Q        Gt  Vt   0��t  �t   0�        uo  1p   S�t  Gu   S�w  Rx   Szz  �z   S�z  �z   S�z  |   S}  �}   S�~  �~   S�  4�   S��  ߀   S��  �   S��  щ   Sj�  ��   S؊  ��   S�  l�   S�  �   S�  $�   Sa�  ��   S        uo  �o   P�t  u   P�w  �w   P�w  x   P�z  �z   P�z  �z   P�~  �~   Pj�  l�   P        �o  �o   P�o  p   W�z  |   W}  �}   W�  4�   W��  �   W��  щ   Wx�  ��   W�  l�   W�  �   W�  $�   Wa�  ��   W        �o  �o   0��z  �z   0��z  {   R{  9{   �T}  9}   0���  �   R�  �   �Tx�  ~�   R~�  ��   �T�  �   R�  $�   0�        {  9{   w#9{  B{   P}  9}   w9}  <}   P�  %�   P        �o  p   P�  �   P�  ��   Q�  $�   P        ��  �   0��  �   0�        �{  �{   P�{  |   �TG�  I�   PI�  ^�   �Ta�  ��   �T        �{  �{   P�{  |   �XR�  T�   PT�  ^�   �Xa�  ��   �X        �{  �{   P�{  �{   t Y�  ^�   P}�  ��   P��  ��   0�        [}  �}   �T��  щ   �T7�  <�   P^�  l�   �T�  �   �T        �}  �}   P�}  �}   Q�}  �}   t ̉  щ   Pg�  l�   P�  ��   Q��  �   �X�  �   P        9}  �}   W��  щ   W�  <�   W^�  l�   W�  �   W        >}  H}   PH}  R}   w�  �   P�  .�   w        u  u   Pu  (u   Q(u  Gu   �T        "x  Rx   P�z  �z   p��z  �z   P        "x  Rx   P        "x  Rx   S        6x  Rx   Q        �~  �~   0��~  �~   Wj�  s�   0�s�  x�   P        ��  ��   P��  ߀   W؊  ��   W        ��  ��   P��  ǀ   Q؊  �   Q�  ��   �T        Pq  Rq   PRq  �q   W�x  y   W�z  �z   W        Yq  \q   P\q  �q   V�x  y   V�z  �z   V        �q  �q   Q�q  �q   t y  y   0��z  �z   P        Zu  mw   S�y  zz   S|  }   S�}  �~   S�~  �~   S4�  b�   S��  ��   S�  _�   S��  ��   S��  s�   S��  ��   Sщ  �   S��  Ȋ   S��  �   Sl�  �   S�  ��   S��  ��   S�  �   S$�  a�   S��  Ԏ   S��  �   S/�  B�   SP�  ��   S��  #�   S        `u  �u   R�u  �u   p �u  �u   s*z  @z   R|  |   R|  %|   p %|  (|   s�|  �|   R�|  �|   p �  �   R~�  ��   R�  ��   Rщ  ԉ   p ԉ  ׉   sP�  V�   R        �u  �u   P�u  v   V��  ��   V͋  �   Vl�  w�   V<�  ��   V^�  ��   VT�  ��   VĐ  ��   V        �u  �u   0���  ��   0���  ބ   Wȅ  �   0�͋  �   Wl�  w�   WT�  k�   0���  ��   W        ��  ބ   v#ބ  �   P��  ��   Pȅ  �   v�  �   P        �u  �u   P�  �   P�  �   Qf�  k�   P        ͋  �   0�l�  w�   0�        (�  *�   P*�  ��   �Tv�  x�   Px�  ��   �TĐ  ��   �T        1�  4�   P4�  ��   W�  ��   P��  ��   WĐ  ̐   Wѐ  ��   W        c�  p�   Pp�  t�   t ��  ��   Pא  ސ   0��  ��   P        ��  ��   �T<�  O�   �Tp�  u�   Pu�  ��   �T^�  ��   �T        H�  K�   PK�  ~�   WJ�  O�   P~�  ��   P^�  |�   W|�  ��   P        �  ��   V<�  ��   V^�  ��   V        �  ��   P��  ��   vO�  R�   PR�  k�   v        Ez  Nz   PNz  uz   W        �|  �|   0��|  }   P�~  �~   p��~  �~   P        �|  }   P        �|  }   S         }  }   W        �  ��   0���  $�   VP�  Y�   0�Y�  ^�   P        ��  �   P�  �   W�  <�   W        �  �   P�  �   V�  <�   V        v  Gv   S�y  �y   S�|  �|   SE~  �~   SK�  [�   S��  ��   S��  ��   S��  Ȋ   S�  �   S        v  Gv   R�y  �y   R�|  �|   R�|  �|   p �|  �|   sE~  R~   RR~  U~   p ��  ��   R��  ��   R��  ��   p ��  ��   s        iv  qv   Pqv  �v   V`�  I�   VN�  n�   V��  ��   V��  D�   V��  ��   V$�  /�   V��  �   V��  �   V�   �   V%�  T�   V��  Đ   V        ^v  �v   0�`�  }�   0���  ��   0���  ֈ   Rֈ  �   �T��  )�   R)�  D�   �T��  ��   R��  ��   �T$�  /�   R��  �   0�        `�  }�   v}�  ��   PN�  d�   P�  �   v#�  �   P        �v  �v   P*�  7�   P7�  ;�   Q�  �   P        ��  D�   0�$�  /�   0�        χ  ч   Pч  N�   �T�  �   P�  ��   �T�  T�   �T        ڇ  ݇   P݇  N�   �X�  �   P�  ��   �X�  T�   �X        �  �   P�  �   t ��  ��   PB�  G�   PM�  T�   0�        &�  ��   �T��  ��   �T֏  ۏ   P��  �   �T��  Đ   �T        ��  ��   P��  ��   Q��  ��   t ��  ��   P�  �   P��  ��   Q��  ��   �X��  Đ   P        �  ��   V��  ۏ   V��  �   V��  Đ   V        	�  �   P�  �   v��  ��   P��  ͏   v        �y  �y   P�y  �y   V        e~  g~   0�g~  �~   PR�  U�   p�U�  [�   P        g~  �~   P        g~  �~   S        {~  �~   V        ��     0�  �   V�  �   0��  �   P        ��  ��   P��  Ê   V�  �   V        ��  ��   P��  ��   Q�  ��   Q��  �   �T        �v  �v   S�y  *z   SL|  �|   S�}  E~   S4�  D�   S��  ��   S��  ��   S��  ͋   S��  #�   S        �v  �v   Q�y  �y   QL|  n|   Q�}  ~   Q4�  :�   Q��  ��   Q��  ��   Q��  ��   Q        w  !w   P!w  mw   �T�  _�   �T��  ~�   �TD�  ��   �Tw�  �   �T/�  a�   �T��  Ԏ   �T/�  B�   �T        w  Hw   0��  �   0��  1�   R1�  c�   �X��  ��   0�D�  n�   Rn�  ��   �Xw�  ��   RQ�  W�   RW�  a�   �X��  Ԏ   0�        A�  c�   �T##c�  l�   P8�  J�   P��  ��   �T#��     P        Ow  Sw   Po�  |�   P|�  ��   Qώ  Ԏ   P        D�  ��   0�w�  ��   0�        ��  ��   P��  8�   �X:�  <�   P<�  Q�   �X��  ��   �X        ��  Â   PÂ  8�   �\E�  G�   PG�  Q�   �\��  ��   �\        �  �   P�  �   t L�  Q�   P��  ��   P��  ��   0�        �  ~�   �X��  ��   �XԌ  ٌ   Pٌ  �   �X/�  B�   �X        A�  D�   PD�  \�   Q\�  `�   t ��  ��   Q��  ��   �\��  ��   P�  �   P=�  B�   P        ��  ~�   �T��  �   �T/�  B�   �T        ǃ  у   Pу  ۃ   �T#��  ��   P��  ˌ   �T#        �y  �y   P�y  z   Qz  *z   �T        ~  ~   0�~  E~   P;�  >�   p�>�  D�   P        ~  E~   P        ~  E~   S        )~  E~   Q        $�  .�   0�=�  A�   QA�  `�   �T��  ��   0���  ��   P        ��  ��   �T        ��  ��   P��  ��   Q��  �   Q�  #�   �X        s  �s   �XGu  Zu   �X�w  �w   P�x  �x   �Xay  �y   �X        [s  ^s   P^s  �s   VUu  Zu   P�x  �x   Pay  y   Vy  �y   P        Rr  �r   t �r  s   �Pmw  �w   t Rx  �x   t �x  �x   �P�x  �x   t �x  �x   t �x  �x   �P�x  �x   t y  ay   t �z  �z   t �~     t   "   �P"  R   t R  a   �Pa  �   t �  
�   �P
�  �   t b�  ��   t ��  ��   �P��  ��   t ߀  ��   t ��  ��   V_�  ��   t ��  ��   �P��  ��   t ��  ��   t ��  ��   �P��  ��   t s�  ��   t ��  ��   �P�  $�   V$�  D�   t D�  j�   VȊ  Ҋ   t Ҋ  ؊   �P��  ��   t ��  ؍   t Ԏ  ގ   t ގ  ��   �P�  /�   VB�  P�   V��  ��   t         Zr  dr   Pdr  �r   t #mw  sw   Psw  �w   t #Rx  bx   t #�x  �x   t #y  y   t #�~  �~   t #�~  �~   t #b�  n�   t #_�  e�   t #        dr  s   SRx  �x   S�x  �x   Sy  ay   S�z  �z   S�~  �   Sb�  ��   S߀  ��   S_�  ��   S��  ��   Ss�  ��   S�  j�   SȊ  ؊   S��  ��   S��  ؍   SԎ  ��   S�  /�   SB�  P�   S��  ��   S        jr  �r   R�r  �r   p �r  �r   sRx  hx   R�x  �x   R�x  �x   p �x  �x   sy  y   Ry  y   p �~  �~   R�~  �~   Rb�  n�   R_�  b�   p b�  e�   s        �r  �r   P�r  s   V  �   V߀  ��   V��  ��   Vs�  ��   V�  j�   VȊ  ؊   V��  ��   V��  ؍   V�  /�   VB�  P�   V��  ��   V        �r  �r   0�  	   0�	  H   W߀  ��   0�s�  ��   WȊ  ؊   W��  ��   0���  ��   W        *  H   v#H  Q   P߀  ��   v��  ��   P��  ��   P        �r  �r   P��  ��   P��  ��   Q��  ��   P        s�  ��   0���  ��   0�        �  �   P�  �   �X/�  1�   P1�  D�   �X��  ؍   �X        �  �   P�  �   W8�  :�   P:�  D�   W��  ؍   W        �  �   P�  �   t ?�  D�   Pƍ  ˍ   Pэ  ؍   0�        �  ��   �X�  $�   �Xe�  j�   P�  /�   �XB�  P�   �X        c�  f�   Pf�  ��   W�  $�   P�  *�   W*�  /�   PK�  P�   P        ��  ��   V�  $�   VD�  j�   V�  /�   VB�  P�   V        �  �   P�  �   vD�  G�   PG�  `�   v        ox  xx   Pxx  �x   �X        -y  /y   0�/y  ay   P�z  �z   p��z  �z   P        /y  ay   P        /y  ay   S        My  ay   Q        b�  q�   0�q�  ��   V        n�  p�   Pp�  ��   WԎ  ��   W        w�  z�   Pz�  ��   VԎ  ��   V        kp  tp   Ptp  }p   V�s  �s   V        �p  �p   R�q  �q   p��q  �q   P        �p  �p   R        �p  �p   S        �p  �p   V        t  t   Pt  Bt   V�w  �w   V        t  "t   P"t  Gt   W�w  �w   W        0�  @�   P@�  f�   Sf�  j�   �P�j�  ��   S��  ��   P��  ƒ   Sƒ  ʒ   �P�ʒ  Ԓ   PԒ  X�   SX�  \�   �P�\�  d�   S        @�  t�   Pt�  ~�   uj�  x�   Px�  |�   u ��  �   P�  �   u \�  b�   Pb�  f�   u m�  z�   PǓ  Փ   PՓ  ؓ   u ��  �   P�  �   u �  �   P�  �   u <�  C�   PC�  F�   u V�  o�   uo�  u�   Pu�  x�   u ��  Ŕ   PŔ  Ȕ   u �  ��   P��  ��   u �  %�   P%�  (�   u L�  T�   PT�  s�   u ��  ��   P��  ��   u �  ��   P��  �   u ;�  B�   PB�  F�   u ��  ��   uǖ  ߖ   u �  �   u9�  Q�   ur�  x�   u~�  ��   u��  ��   uݗ  ��   u�  .�   uO�  _�   ue�  }�   u8�  >�   u g�  q�   u        `�  e�   P        ^�  t�   1�t�  Y�   0�Y�  b�   1���  <�   1�<�  o�   0�o�  ��   1���  3�   1�3�  ;�   0�;�  ��   1���  ՗   0�՗  ݗ   1�ݗ  �   0��  g�   1�g�  s�   0�s�  C�   1�C�  ��   0���  Л   1�Л  �   0��  6�   1�6�  ��   0���  ��   1���  Ǟ   0�Ǟ  �   1��  �   0��  v�   1�v�  �   0��  |�   1�|�  ��   0���  ʢ   1�ʢ  ڢ   0�ڢ  �   1��  ��   0���  ��   1���  �   0��  �   1��  ��   0���  �   1��   �   0� �  C�   1�C�  d�   0�        t�  Y�   SC�  ��   SЛ  �   S6�  ��   S��  Ǟ   S�  �   Sv�  �   S|�  ��   Sʢ  ڢ   S�  ��   S��  �   S�  ��   S�   �   SC�  d�   S        w�  Y�   WC�  ��   WЛ  �   W6�  ��   W��  Ǟ   W�  �   Wv�  �   W|�  ��   Wʢ  ڢ   W�  ��   W��  �   W�  ��   W�   �   WC�  d�   W        ~�  Y�   SC�  ��   SЛ  �   S6�  ��   S��  Ǟ   S�  �   Sv�  �   S|�  ��   Sʢ  ڢ   S�  ��   S��  �   S�  ��   S�   �   SC�  d�   S        ��  ˑ   Pˑ  ё   uC�  U�   PЛ  ԛ   Pԛ  �   u6�  C�   PC�  F�   uv�  ��   P��  ��   P��  ��   u��  ��   P��  ��   u|�  ��   u�  �   P�  ��   u        ֑  ޑ   Pޑ  #�   V�  �   VȠ  �   Vʢ  ڢ   V�  ��   V��  �   V�   �   V        ˑ  �   0��  �   0��  .�   UȠ  �   0���  �   Uʢ  ڢ   U��  ţ   0��   �   U        �  .�   v#.�  ?�   PȠ  �   v�  �   P��  ��   P        �  �   Pء  �   P�  �   Q��  ţ   P        ��  �   0��   �   0�        u�  w�   Pw�  �   �H�  L�   �HУ  ң   Pң  �   �H        ~�  ��   P��  �   U�  L�   U٣  ۣ   Pۣ  �   U        ��  ��   P��  ��   t :�  ?�   PE�  L�   0��  �   P        ��  ��   �H�  �   �Hm�  r�   Pr�  ��   �H        L�  O�   PO�  ��   U��  ��   P��  �   U�  �   P{�  ��   P        �  ��   V�  �   VL�  ��   V        �  ��   P��  ��   vL�  O�   PO�  h�   v        Z�  v�   Pv�  z�   Qz�  ��   �H        X�  ��   R��  ��   p���  ��   P        X�  ��   R        X�  ��   S        j�  ��   P        v�  ��   0���  ��   V�  ��   0���  ��   P        ��  ��   P��  ��   VC�  d�   V        ��  ��   P��  ��   UC�  d�   U        ��  ��   P��  ǒ   Vʒ  ��   V        ��  ʒ   R        ��  ƒ   Sƒ  ʒ   �P�        �  ��   W        Y�  b�   �\0�  Q�   PQ�  T�   s 2$q "T�  \�   r2$q "        Y�  b�   S0�  X�   SX�  \�   �P�        \�  m�   S        m�  ��   S�  8�   SY�  �   Ss�  C�   S  Л   S�  6�   S��  ��   SǞ  �   S�  v�   S�  |�   S��  ʢ   Sڢ  �   S��  ��   S�  �   S��  �   S �  C�   S        z�  ��   P��  ��   r ��  ��   p ��  ��   v ��  ��   W�  �   PY�  c�   r         ��  ��   P��  ��   W�  8�   W        Y�  �   Ss�  C�   S  Л   S�  6�   S��  ��   SǞ  �   S�  v�   S�  |�   S��  ʢ   Sڢ  �   S��  ��   S�  �   S��  �   S �  C�   S        \�  �   Vs�  C�   V  Л   V�  6�   V��  ��   VǞ  �   V�  v�   V�  |�   V��  ʢ   Vڢ  �   V��  ��   V�  �   V��  �   V �  C�   V        c�  �   Ss�  C�   S  Л   S�  6�   S��  ��   SǞ  �   S�  v�   S�  |�   S��  ʢ   Sڢ  �   S��  ��   S�  �   S��  �   S �  C�   S        g�  ��   P��  ��   us�  ��   P��  ��   P��  Ě   u�  ��   P��   �   u  ě   Pě  ț   u(�  *�   P*�  .�   um�  w�   P�  ��   u��  ��   P��  ¢   u        ��  Ù   PÙ  �   W��  h�   W��  ��   W��  ��   W0�  v�   W�  "�   WC�  |�   Wڢ  �   W��  ��   W�  �   W��  �   W �  C�   W        ��  �   0���  ��   0���  ��   0���  �   U0�  v�   U�  "�   U�  �   U��  �   0�        ��  ��   w��  ��   Pɝ  �   w#�  �   P��  ��   P        �  ��   P\�  i�   Pi�  m�   Q�  �   P        0�  v�   0��  �   0�        �  ��   P��  m�   �H��  ��   P��  �   �H��  ��   �H        ��  ��   P��  m�   U�  �   P�  �   U��  ��   U        -�  :�   P:�  >�   t �  �   P��  ��   P��  ��   0�        �  ��   �Hd�  i�   Pi�  |�   �Hڢ  �   �H �  C�   �H        N�  Q�   PQ�  ��   Uw�  |�   P�  �   P �  >�   U>�  C�   P        �  ��   WC�  |�   Wڢ  �   W �  C�   W        �  ��   P��  ��   wC�  F�   PF�  _�   w        ��  ��   PǞ  ɞ   Pɞ  �   W        �  C�   P�  �   p��  �   P        �  C�   P        �  C�   S        $�  C�   W        m�  w�   0�w�  ��   W��  Ţ   0�Ţ  ʢ   P        ��  �   P�  +�   W"�  C�   W        �  �   P�  0�   U"�  C�   U        o�  ��   S        ��  ��   P��  ��   V        ��  ��   P��  ��   t         T�  c�   Pc�  s�   u8�  >�   u        8�  Y�   S        ;�  K�   P��     P        �  &�   V��&�  )�   V�U��)�  -�   V�U�W��-�  0�   V�U�W�P��0�  4�   V�U�W�s(��4�  6�   V�U�W�s(�P�6�  :�   V�U�W�s(�s0�:�  g�   V�U�W��H��L���  ��   V�U�W��H��L���     �U�W��H��L�        �  g�   � �  ��     � �          �  g�   S��     S        G�  g�   � �          G�  g�   S        ��     Q        ��     S        �  ;�   V        �  ;�   S        �  ;�   P        b�  ��   P��  ��   s 2$q "��  ��   r2$q "        b�  ��   S        ��  ��   l4	���     p  ǖ   l4	�        ��  ǖ   S        ��  ǖ   P        ǖ  ��   D4	���  ��   p��   �   D4	�        ǖ   �   S        �   �   P         �  0�   4	�0�  4�   p4�  9�   4	�         �  9�   S        �  9�   P        9�  i�   04	�i�  m�   pm�  r�   04	�        9�  r�   S        T�  r�   P        ~�  ��   X4	���  ��   p��  ��   X4	�        ~�  ��   S        ��  ��   P        ݗ  �   �4	��  �   p�  �   �4	�        ݗ  �   S        ��  �   P        �  F�   4	�F�  J�   pJ�  O�   4	�        �  O�   S        1�  O�   P        e�  �   Sg�  s�   S        ��  ��   R        p�  ��   P��  	�   S	�  �   �P��  O�   S        ��  ��   �\���  	�   V�  O�   V        ��  ��   P��  ¤   Q�  	�   P        ��  ��   R֤  �   R�  +�   R        P�  Z�   PZ�  ��   S��  ��   �P���  ��   S        P�  e�   R��  ��   R        e�  ��   V��  ��   P��  ��   V        l�  }�   P}�  ��   t         Z�  e�   p ��  ��   p ��  ��   s        ��  ʥ   Pʥ  ˥   �P�˥  �   P�  	�   S	�  
�   �P�
�  �   S�  �   �P�        �  ��   P��  ��   R��  �   P
�  �   P         �  .�   P.�  G�   �\G�  ��   S��  ֧   �\        H�  ��   W>�  G�   WG�  ^�   R^�  ��   W        e�  n�   Pn�  x�   �\#1x�  ��   �[G�  `�   P`�  k�   s1k�  ��   �[        y�  ��   P��  ��   r        y�  ��   �[�H$H&0���  ��   qP���  ��   Q        y�  ��   �\        ��  ��   R        ��  ��   P��  ��   r        ��  ��   �[�H$H&0���  ��   qP���  ��   Q        Ԧ  4�   R��  ��   R        Ԧ  4�   �T��  ֧   �T        Ԧ  �   P�  4�   P��  ��   P��  ��   �Tr O%�T"r 1&r "�        Ԧ  �   U�  4�   U��  է   Uէ  ֧   p        ��  է   Uէ  ֧   p        r�  ~�   P~�  ��   Q        c�  ��   V        �  �   P�  ��   S��  ��   �P���  6�   S6�  :�   �P�:�  ݫ   S        ��  ��   P��  ��   U��  �   P�  �   P�  "�   U:�  P�   PP�  ��   U��  ��   P        �  )�   R)�  C�   p ��  ��   R�  ��   R�  �   p ��  ܩ   R�  �   R��  ��   R��  ��   p ˫  ҫ   Rҫ  ի   p         ;�  ��   S        Y�  ��   P��  ��   u        a�  ��   S        x�  ��   U        �  ��   U        �  ��   S        ��  �   U�  �   P        ��  �   B��  �   r         ͨ  ڨ   Pڨ  ި   t         �  ��   S        5�  L�   PL�  ��   W        T�  ��   P��  ��   u        \�  ��   S        w�  ��   U        ��  ��   U        ��  ��   S        ��  �   S��  ݫ   S        ��  �   Q�  �   u�  �   5��  �   3�%�  ,�   4�        Ū  �   �\�  ��   V        Ū  �   Q�  �   u        Ū  �   S        ڪ  �   U        ڪ  �   �\�  ��   V        ڪ  �   Q�  �   u        O�  ��   Q��  ��   u��  ��   5���  ��   4���  ��   3�        [�  |�   �\|�  ��   W        [�  ��   Q��  ��   u        [�  ��   S        m�  ��   U        m�  |�   �\|�  ��   W        m�  ��   Q��  ��   u        �  �   P�  .�   V.�  1�   �P�1�  P�   VP�  S�   �P�S�  ��   V��  ��   P��  Ԯ   VԮ  �   P�  ��   V��  ��   �P���  ��   V        �  �   p �  �   R�  �   v1�  F�   RS�  p�   Rp�  x�   v.�  6�   Rt�  ��   R��  ��   p ��  ��   v­  ܭ   R        7�  P�   PP�  t�   S��  ��   P��  ��   W��  ��   S��  ��   Q��  ��   S��  ­   P�  �   P�  >�   W        �  %�   VL�  ��   V��  ��   �P���  k�   V        �  %�   PL�  S�   PS�  ��   S��  !�   S&�  7�   S<�  k�   S        q�  u�   Pu�  ��   Wӯ  ׯ   Pׯ  �   R�  �   R�  &�   �L&�  <�   W        b�  ��   	����  ¯   	��¯  ʯ   Pʯ  &�   U&�  <�   	��        �  �   R        �  �   U        �  �   V        ��  �   W        i�  .�   V>�  ��   V��  ��   P��  Ԯ   VԮ  �   P�  L�   Vk�  ��   V        ��  ��   P��  .�   U>�  L�   Uk�  ��   U        ��  ��   P��  .�   �L>�  L�   �Lk�  ��   �L        ��  .�   V>�  ��   V��  ��   P��  Ԯ   VԮ  �   P�  L�   Vk�  ��   V        ��  ��   0���  .�   W>�  ��   W��  ��   P��  Ү   WԮ  )�   W1�  L�   Wk�  ��   W        ��  ��   S�  �   S��  ��   SԮ  �   S        ��  ��   1�G�  T�   1�T�  `�   R��  ��   1�ʮ  �   1���  	�   4��  1�   1�        G�  \�   P\�  `�   t ��  ��   Pʮ  Ԯ   P�  �   P��  	�   P�  1�   PG�  L�   P        s�  ��   W        s�  ��   V        ��  ��   rԮ  �   r        E�  P�   PP�  t�   S        E�  t�   V        ��  ��   1��  >�   0�        �  >�   W        �  >�   V        ��  ��   P��  f�   Sf�  j�   �P�j�  ��   S��  ��   �P���  �   S�  �   �P��  Զ   S        ��  ٰ   Rٰ  h�   Wh�  j�   �R�j�  v�   Rv�  ��   �R���  ��   W��  �   �R��  �   W�  O�   �R�O�  g�   Wg�  Զ   �R�        ��  ٰ   Qj�  s�   Qs�  y�   p         հ  ٰ   Rٰ  h�   Wh�  j�   �R���  ��   W�  �   W�  �   �R�O�  g�   W        հ  f�   Sf�  j�   �P���  ��   S�  �   S�  �   �P�O�  g�   S        �  ��   P��  -�   s��  ��   s�  ��   sO�  g�   s        ް  �   P�  g�   Vg�  j�   P��  ��   V�  �   VO�  g�   V        ��  ��   P        E�  `�   R        j�  ��   S��  ��   �P���  �   S�  O�   Sg�  Զ   S        g�  L�   S@�  ��   S��  Զ   S        g�  ��   0���   �   �\ �  +�   P+�  D�   �\D�  L�   P@�  ��   �\��  Զ   �\        g�  ��   0��  �   P�  �   t ��  ��   P        x�  ��   P��  ��   U        ��  ��   0���  Ʋ   0�Ʋ  ��   V��  L�   0�@�  ��   2���  ��   0���  Զ   2�        ��  Ʋ   PƲ  �   w @�  D�   PD�  T�   w T�  Y�   $���  ˶   w         ��  �   W��  L�   W@�  z�   W��  ��   W��  Զ   W        Y�  ��   Q˶  Զ   Q        Y�  ��   S˶  Զ   S        p�  ��   P        ��  ��   P��  ��   V        ��  ��   P��  �   V        ��  Ĵ   P        ̴  ݴ   Pݴ  �   Q        �  �   P�  =�   S=�  A�   �P�A�  ̷   S̷  ٷ   Pٷ  '�   S'�  4�   P4�  ��   S��  ��   �P���  Ź   SŹ  ۹   P۹  ܹ   �P�ܹ  �   P�  �   �P��  �   S        �   �   RA�  u�   R̷  �   R'�  P�   R_�  j�   R��  ۹   Rܹ  �   R�  �   R@�  M�   R�  ��   R	�  �   R        !�  7�   Pú  Һ   PҺ  �   V        z�  ��   P��  ̷   Un�  _�   U�  ú   UM�  �   U�  ~�   U��  	�   U        o�  ��   0�n�  z�   0�z�  ��   R��  ��   R�  �   0�u�  ��   0���  ��   R��  	�   R        ��  ��   �X#��  ĸ   P�  �   u�  3�   PM�  f�   P�  �   P        ��  ��   P��  ��   P��  Ȼ   PȻ  ̻   Q        ��  ջ   0���  	�   0�        �  _�   �X.�  C�   �Xy�  ~�   P��  ��   �X��  ݼ   �X        $�  '�   P'�  Z�   V>�  C�   P��  ��   P��  ؼ   Vؼ  ݼ   P        ��  _�   U.�  ~�   U��  ��   U��  ݼ   U        Ƹ  и   Pи  ڸ   uC�  S�   PS�  p�   u        M�  O�   PO�  ��   V�  �   P�  .�   V��  ��   Vݼ  ��   V        Y�  \�   P\�  ú   W"�  $�   P$�  .�   W��  ��   Wݼ  ��   W        ��  ��   P��  ��   t )�  .�   P��  ��   0���  ��   P        �  �   p��  '�   PH�  M�   0�        ��  '�   P        ��  '�   S        �  '�   V        _�  j�   0�j�  ��   W�  ��   0���  �   P        �  �   P�  ;�   V~�  ��   V        �  (�   P(�  @�   W~�  ��   P��  ��   W         �  T�   P��  �   P         �  7�   R7�  ̿   u�|̿  d�   ��|         �  K�   QK�  ̿   u�|̿  ��   ��|��  �   Q�  d�   ��|        ��  ��   V�  �   V!�  .�   V<�  f�   VG�  d�   V        ��  ��   P��  ʿ   V�  !�   0�.�  4�   P4�  <�   V        �  !�   P        ��  {�   u�|�{�  о   Wо  ̿   u�|�̿  Ϳ   ��|��  '�   ��|�'�  +�   P+�  H�   ��|�H�  G�   WG�  M�   ��|�M�  d�   W        ��  Ľ   PĽ  ��   u�}�  �   ��}!�  +�   ��}<�  \�   ��}G�  ^�   ��}        ��  Ϳ   A��  d�   A�        ��  ��   S��  Ϳ   �P��  �   S�  !�   �P�!�  K�   SK�  \�   w \�  h�   s~�h�  G�   �P�G�  P�   SP�  ^�   w ^�  d�   ss�        3�  ��   q �  �   q !�  +�   q <�  \�   q G�  ^�   q         5�  u�   t u�  ��   u�}��  ��   t��  ��   t �  �   t !�  h�   t v�  ��   t G�  d�   t         f�  ��   R��  ��   u�|��  о   �P#�G�  R�   RR�  X�   ��|X�  ^�   w #�^�  d�   s~�        f�  {�   u�|�{�  о   WG�  M�   ��|�M�  d�   W        �  Ϳ   A�        �  ̿   u�|̿  Ϳ   ��|        �  ̿   u�|̿  Ϳ   ��|        �  ʿ   V        �  �   u�}��  ɿ   Sɿ  ̿   u�}�̿  Ϳ   ��}�        ��  ��   r ��  ��   t ��  ��   uL        ��  ��   t         ��  ɿ   Sɿ  ̿   u�}�̿  Ϳ   ��}�        �  �   1�<�  G�   1�        �  �   ��|�<�  H�   ��|�H�  G�   W        f�  h�   Ph�  v�   Vv�  �   P�  �   V�  �   P�  G�   V         �  G�   V         �  G�   W         �  G�   R        ��  ��   S��  ��   Q��   �   S �  '�   R'�  G�   S        ��   �   P �  �   t         *�  ��   u�}1��  �   ��|1�!�  +�   ��|1�<�  \�   ��|1�G�  ^�   ��|1�        b�  v�   p�v�  ��   uT1�        ��  ��   q���  ��   u`1�        .�  C�   WC�  E�   P��  ��   W        ��  D�   UE�  Y�   Ui�  ��   U��  ��   0���  ��   U        ��  _�   A�i�  ��   A�        ��  _�   �ܥ  i�  ��   �ܥ          ��  ��   P��  _�   � i�  ��   �         ��  
�   PE�  Y�   P��  ��   P��  ��   P��  ��   P        ��  _�   0�i�  ��   0�        ��  �   T�  �   �P��  �   T�  1�   �P�1�  >�   T>�  E�   �P�E�  _�   Ti�  s�   Ts�  ��   �P���  ��   T��  ��   �P���  ��   T        ��  �   P           8    Q�R�8   H    Q���H   Q    ����Q   �    P�R��   �    P����   �    �����   �    P�R��   �    Q�R��   �    Q����   �    P�R��   �    P����      Q���     P�R�  +   Q�R�+  9   ����        #   8    Q�R�<   @    Q�R�H   J    Q�R�~   �    P�R��   �    Q�R�  +   Q�R�        !   <    Q<   H    UQ   q    Pq   �    �l�   �    P�   �    Q�   �    P�      Q     P  +   Q        !   8    R8   H    �Q   q    Rq   �    �h�   �    R�   �    ��   �    R�      �  +   R        !   D    � Q   �    � �   �    � v $��   �   + � O�(  / 0@K$(	 1$#/���O'$��   �    �   !   � +  4   � v $�4  9  + � O�(  / 0@K$(	 1$#/���O'$�        !   D    �D   H    RQ   �    ��   �    W�   �    R�   �    U�   !   �+  9   U        �   �    R�   �   
 t q �%�        �   �    P�   �    W�   �    w��   �    P!  +   1�+  9   W        D   F    PF   H    V�   �    0�        q   |     v �|   �    U�   �     v ��   �   *  O�(  / 0@K$(	 1$#/���O'�+  4    v �4  9  *  O�(  / 0@K$(	 1$#/���O'�        h   k    v O'�k   �    V�   �   ' O�(  / 0@K$(	 1$#/���O'�  4   V4  9  ' O�(  / 0@K$(	 1$#/���O'�        �   �    R�   �    t +  9   t         �   �    P+  2   P        @   G    P�R�|   �    P�R��   �    P�R�X  _   P�R�           8    W�P�8   :    W�R�:   E    W���E   G    ����G   x    W�P�x   |    W�R�|   �    W����   �    �����   �    W�P��   �    W�R��   �    W����   �    W�P��   �    W�R��   �    W����   �    �����   �    W�P��   �    W�R��   �    W����   _   ����_  u   W�P�               Q�P�   D    Q�V�D   G    Q���G   t    Q�V�t   �    � ����   �    Q�V��   �    Q����   �    Q�V��   �    � �V��   _   � ���_  d   Q�V�d  h   Q���h  u   � ���        0   <    WG   �    W�   �    ��   �    W�   �    U�   �    W�   �    ��   �    �\_  u   W        0   8    P8   :    R:   G    �G   x    Px   |    R|   �    ��   �    P�   �    R�   �    ��   �    P�   �    R�   �    ��   �    �`_  u   P        0   <    QG   t    Q�   �    Q�   �    Q�      �   #   V#  G   �dG  I   P_  h   Qh  p   �         0   <    VG   t    V�   �    V�   �    R�   �    V�   �    ��   �    V�   	   �	     P     v �h��%�q �$!�     �l�h��%�q �$!�     �l�h��%�u �$!�  ?   Q?  X   R_  d   Vd  p   �        �   �    P�   !   W!  _   ��h��%�        �   �    0�_  u   1�        t   |    0��   �    0�;  X   0�        �   �     u ��   �    P�   �    W�      R  _   �h        W   Z    u O'�Z   `    U`   x   & Op (  / 0@K$(	 1$#/���O'�x   |   & Or (  / 0@K$(	 1$#/���O'�|   �   ' O�(  / 0@K$(	 1$#/���O'��   ^   U^  _  ' O�(  / 0@K$(	 1$#/���O'�_  u  & Op (  / 0@K$(	 1$#/���O'�        !  ;   R;  P   W        !  ;   P;  \   V                P   A    P            	    R	   @    U@   A    �R�            	    0�	   !    Q!   #    qy�#   A    Q           /    R/   =    p            	    0�	   ?    W?   @    u @   A    �R        P   �    P�   �    V�   �    P�      W  8   P@  G   WG  Y   �LY  c   r�c  y   r�y  �   R�  �   P�  �   W�  �   �L�  �   W�  �   �L�  �   W�     v�     v�     V  $   P$  '   W'  �   �L�  �   W�  �   �L�  �   P�  �   W�  �   �L�  �   P�  �   W�  �   �L�  �   P�  �   W�     r�     r�  &   p�&  3   v�3  I   v�I  Q   VQ  r   Pr  {   W{  �   v��  �   v��  �   V�  �   W�  �   v��  �   v��  �   V�  �   W�     v�     v�  %   V%  2   P2  ;   W;  C   v�C  ]   v�]  b   p�b  s   r�s  �   r��  �   P�  �   W�  �   �L�  �   W�     �L     W     r�  0   r�0  <   w�<  C   v�C  Y   v�Y  s   Vs  |   W|  �   v��  �   v��  �   V�  �   P�  �   W�  �   v��  �   v��  �   V�  �   P�  �   W�     �L     r�  -   r�-  2   P2  9   W9  C   r�C  _   r�_  s   Rs  w   �Lw  �   r��  �   R�  �   r��  �   P�  �   W�  �   r��  �   r��  �   p��  �   P�     W     r�  1   r�1  ;   p�<  ^   P^  i   Wi  �   P�  �   W�  �   r��  �   r��  �   p��  �   v��  �   v��  �   V�     P  	   W	     r�  .   r�.  2   p�3  Z   PZ  a   Wa  s   r�s  �   r��  �   R�  �   �L�  �   r��  �   R�  �   r��  �   P�  �   W�  �   �L�   	   P	  E	   PE	  j	   �Lx	  +
   �L        P   �    R�   �    �D�   +
   �R�        P   �    �         P   �    �        S   �    0��   8   ��@  �   ���  k   ��r  �   ���  �   p��  �   ���     P  �   ���  �   ��  S   ��Z  @	   ��E	  +
   ��        �   �    �         �   �    R�   �    p �   �    R�   �    p �      w@  E   RE  J   VJ  N   p N  �   �L1�  �   R�  �   p �  �   w�  �   �L1�  �   w�  �   p �  �   p �     �L1$  �   p �  �   p~�  �   p �  �   p}�  �   p �  �   p{�  �   p �      �L1r  {   p {  �   �L1�  �   p �  �   �L1�  �   p �  -   �L12  ;   p ;  `   �L1�  �   p �  �   �L1�  �   p �  �   w�  �   �L1     p   8   �L1s  |   p |  �   �L1�  �   p �  �   �L1�  �   p �  �   �L12  9   p 9  _   �L1�  �   p �  �   �L1�     p   7   �L1^  d   p d  h   w�  �   p �  �   �L1  	   p 	  2   �L1Z  a   p a  �   �L1�  �   p �  �   w�  �   �L1E	  K	   p x	  ~	   p ~	  �	   pw�	  �	   p �	  �	   p}�	  �	   p �	  �	   �L1�	  �	   p �	  �	   �L1�	  �	   p �	  �	   p}�	  �	   p �	  �	   �L1�	  
   p 
  +
   �L1        T  V   PV  �   �@�  �   Q�  �   P�  �   r ��  $   V$  X   �LX  r   V�  �   W�  �   W  2   WW  b   Wb  �   �L�  �   R�  �   �L_  u   V�  �   V�  �   V�  �   �L�     V)  Z   V�  �   V�   	   W 	  @	   �L@	  E	   V        y  �   W  $   WI  N   WN  X   R)  :   V:  <   p�<  Y   �#�Y  \   W\  s   R�  �   W�  �   W)  2   V�  �   V)  ?   V�  �   W�  �   R�  �   V	  #	   W        �  �   WX  r   R�  �   R�     R@  Z   R#	  4	   W4	  E	   w �        T  �   �S�          T  Y   �LY  c   r�c  �   r��  �   p�        T  Y   0�Y  q   Qq  s   qy�s  �   Q        g  }   V}  �   P�  �   r�  �   p        T  Y   0�Y  �   W        �  �   ���  .  �   ���  E	  
   ���          �  �   �L.  �   �LE	  
   �L        �  �   W.  u   Wu  �   QE	  K	   Qx	  �	   Q�	  �	   W�	  �	   Q�	  �	   W�	  �	   �#��	  �	   Q�	  �	   W�	  �	   Q�	  
   W        �  �   � .  �   � E	  
   �         a  j   �         �	  
   �         
  
   �         j  �   ���  E	  �	   ���  �	  �	   ���  
  
   ���          j  �   �LE	  K	   �LK	  x	   Px	  ~	   �L~	  �	   P�	  �	   �L�	  �	   P�	  �	   �L�	  �	   P�	  �	   �L�	  �	   P�	  �	   �L�	  �	   P
  
   P        j  �   �@E	  �	   �@�	  �	   �@
  
   �@        j  u   Wu  �   QE	  K	   Qx	  �	   Q�	  �	   Q�	  �	   W�	  �	   �#��	  �	   Q�	  �	   W�	  �	   Q�	  �	   W        j  �   �LE	  �	   �L�	  �	   �L
  
   �L        H	  j	   R{	  �	   R�	  �	   R�	  �	   R�	  �	   R�	  �	   r 
  
   r         �	  �	   P        �	  �	   Q�	  �	   qy��	  �	   Q        �	  �	   R�	  �	   p        �	  �	   W�	  �	   R        �	  �	   �L�	  �	   R        �     v�     v�  $   p�        �     Q     qy�  $   Q          $   R        �  $   W        �     r�     r�  &   p�&  3   v�3  Q   v�Q  r   p�        �     Q     qy�  "   Q          &   W        �  $   V$  k   �L          r   �S�               r�  &   p�&  3   v�3  Q   v�Q  r   p�          &   0�&  A   QA  C   qy�C  d   Q        7  I   RI  Q   vQ  k   p          &   0�&  N   WN  X   R        {  �   v��  �   v�        {  �   Q�  �   qy��  �   Q        �  �   R        {  �   W        �  �   v��  �   v�        �  �   Q�  �   qy��  �   Q        �  �   R        �  �   W        �     v�  %   v�%  2   p�        �     Q     qy�  2   Q          2   R        �  2   W        �  �   V        ;  C   v�C  ]   v�]  b   p�b  s   r�s  �   r��  �   p�        ;  Q   QQ  S   qy�S  [   Q        G  b   R        ;  b   Wb  �   �L        W  �   �4�          W  ]   v�]  b   p�b  s   r�s  �   r��  �   p�        W  b   0�b  �   Q�  �   qy��  �   Q        w  �   W        W  b   0�b  �   V        �  �   P�  �   w�&
  +
   P        �     P     ��             r�  0   r�0  <   w�<  C   v�C  s   v�          !   Q!  #   qy�#  2   Q          .   W.  0   r0  8   w          :   V:  <   p�<  s   �#�        8  s   �S�          8  <   w�<  C   v�C  s   v�        8  <   0�<  Q   QQ  S   qy�S  s   Q        G  Y   RY  d   v        8  <   0�<  \   W\  s   R        |  �   v��  �   v��  �   p�        |  �   Q�  �   qy��  �   Q        �  �   R        |  �   W        �  �   v��  �   v��  �   p�        �  �   Q�  �   qy��  �   Q        �  �   R        �  �   W          2   �S�               �L     r�  2   r�             0�  !   Q!  #   qy�#  2   Q          2   W             0�  2   V        9  C   r�C  s   r�s  w   �L#�w  �   r��  �   r�        9  Q   QQ  S   qy�S  w   Q        G  w   W        9  u   V        p  �   �S�          p  s   Rs  w   �Lw  �   r��  �   r�        p  w   0�w  �   Q�  �   qy��  �   Q        �  �   W        p  w   0�w  �   V        �  �   r��  �   r��  �   p�        �  �   Q�  �   qy��  �   Q        �  �   W        �  �   V             r�  1   r�1  ;   p�          !   Q!  #   qy�#  ;   Q          ,   W,  .   P.  1   r1  7   p          ?   V        �  �   r��  �   r��  �   p��  �   v��  �   v��     p�        �  �   Q�  �   qy��  �   Q        �  �   W        �  �   V�  �   �L        �     �S�          �  �   r��  �   p��  �   v��  �   v��     p�        �  �   0��  �   Q�  �   qy��  �   Q        �  �   R�  �   v�  �   p        �  �   0��  �   W�  �   R        	     r�  .   r�.  2   p�        	  !   Q!  #   qy�#  2   Q          6   W        	  Z   V        a  s   r�s  �   r��  �   �L#��  �   r��  �   r�        a  �   Q�  �   qy��  �   Q        w  �   W        a  �   V        �  �   �S�          �  �   R�  �   �L�  �   r��  �   r�        �  �   0��  �   Q�  �   qy��  �   Q        �  �   W        �  �   0��  �   V        �   	   P        �  �   Q�  �   qy��  �   Q        �   	   V        �   	   W 	  @	   �L        �  E	   �S�          �  E	   P        �   	   0� 	  	   Q	  	   qy�	  2	   Q        	  	   V	  7	   R7	  >	   p        �   	   0� 	  #	   W        0
  @
   P@
  �
   V�
  �   ���  �   V�  �   �P��  �   ��        0
  �
   R�
  �   U�  �   �R��  �   U        �
  �
   P�
  �
   Q�
  �   ���  �   ��        �
  �
   P�
  �
   W�
  �   ���  �   ���  V   ���  �   W�  &   ���     ��  �   ��        �     ��#�  ,   VG  \   V�  �   ��#�Y  �   V�     V�  �   ��#�          P   0�P  \   W^  �   W�     0�        �  �   ����"#��  �  
 ��r "#��  �   R^  h   ����"#�h  p  
 ��p "#�p  v   R        �
  �
   V�
  �   ���  �   ��        �
  �   U�  �   U        �
  �
   P�
  �
   V�
  �   ���  �   w��  �   W�  �   w��  �   W�     ��  ,   w�,  .   W.  �   w��  *   w��  �   V�  �   W�  9   ��9  <   w�<  H   WH  \   w�f  v   w��  �   W�  �   w��     �L1�  &   w��  	   w�  p   w�p  �   ���  �   w�        �
     P)  9   P<  @   P@  V   Vw  �   V�  �   V�  �   v��  �   V�     v�     V  &   v�&  �   V�     V�  �   P�     V'  \   Vf  v   Vv  �   �D1��  �   V�  �   �D1��  �   V�  �   V�  �   �D1��  �   V�     �D1�     V     �D1�  !   V!  &   �D1�  I   VI  P   �D1�P  p   Vp  �   P�  �   V�  �   V�  �   V        �
  �   0��  �   ���     0�  �   ���  j   ���  9   0�9  ?   P?  \   ��f  &   ���  p   ��p  �   0��  �   ��        )  <   Vw  }   W'  .   W          9   P          !   Q!  #   qy�#  9   Q          5   W          <   V        V  }   V        V  q   Qq  s   qy�s  }   Q        g  }   R        V  }   W        9  �   �4�  f  �   �4�  �  &   �4�    p   �4�          9  �   v�f  v   v�v  �   �D�  �   v��  �   �D�  �   v��  �   �D�  �   v��     �D     v�     �D  !   v�!  &   �D  I   v�I  P   �DP  p   v�        9  >   P>  �   ��f  �   ���  &   ��  p   ��        9  �   ��f  �   ���  &   ��  p   ��        �  �   �4�  f  �   �4�  �  &   �4�  9  P   �4�          �  �   v�f  v   v�v  �   V�  �   v��  �   V�  �   v��  �   V�  �   v��     �D     v�     P  !   v�!  &   V9  I   v�I  P   V        �  �   �Hf  �   �H�  &   �H9  P   �H        �  �   ��f  �   ���  &   ��9  P   ��        �  �   v�f  v   v�v  �   �D�  �   v��  �   �D�  �   v��  �   �D�  �   v��     �D     v�     �D  !   v�!  &   �D9  I   v�I  P   �D        s  �   R�  �   P�  �   p �  �   R�  �   R     R  &   RF  K   p K  P   P        �     V        �  �   Q�  �   qy��     Q        �  �   R�     v        �  �   W�     R        F  K   PK  P   v|�        i  t   ��        P  `   ��        `  p   ��        �  �   P�  �   p|�          H   V          !   Q!  #   qy�#  H   Q          H   R          .   W        �
  �
   Q�
  �   ���  �   ��        �  �   ��  \  �   ��  &  Y   ��  �  �   ��  �  �   ��          �  �   V\  �   V&  -   V�  �   V�  �   ���  �   V�  �   V�  �   v}��  �   V        �  �   ��\  �   ��&  Y   ���  �   ���  �   ��        �  �   ��\  �   ��&  Y   ���  �   ���  �   ��        �  �   ��        �  �   ��        �  �   ��        �  �   ��  &  Y   ��  �  �   ��  �  �   ��          �  �   V&  -   V-  Y   R�  �   V�  �   R�  �   V�  �   ���  �   V�  �   R�  �   V�  �   P�  �   R�  �   V�  �   R�  �   V�  �   v}��  �   R        �  �   ��&  Y   ���  �   ���  �   ��        �  �   ��&  Y   ���  �   ���  �   ��        �  �   V&  -   V�  �   V�  �   ���  �   V�  �   V�  �   v}�        -  A   QA  H   PH  J   p �  �   P�  �   P�  �   P�  �   P�  �   v         �  �   R        �  �   Q�  �   qy��  �   Q        �  �   V�  �   P        �  �   W�  �   Q        �  �   V�  �   v}��  �   V        �  V   ���  �   ���     ���  �   ��        �  �   u��  �   P�  �   u��  �   u�&  -   u��  �   u��     u��  �   u��  �   P�  �   u�        G  P   W        ,  \   V        ,  A   QA  C   qy�C  \   Q        7  \   R        ,  P   W        ^  �   ��        �     P  ,   U,  6   P6  j   Wj  �   P�  �   W�  �   P�  �   W�     W      P   +   W+  0   P0  ;   W;  @   P@  K   WK  P   PP  �   W�  "   p�"  4   W4  C   w�C  �   W�  �   P�  +   W+  I   RI  X   p�X  ]   P]  ~   W~  �   P�  K   WK  O   PX  f   W�  �   W�  �   w��  �   W�      P   :   W:  S   p�S  �   ��}1��  �   W�  �   P�  �   p��  �   ��}1��  �   W�     p�     v�     ��}1�  '   p�'  7   W7  b   Rb  >   W>  B   p�B  T   ��}1�T  [   p�[  `   ��}1�`  g   p�g  l   ��}1�l  p   p�p  �   ��}1��  �   R        �  ,   R,  �   ��}          ,   1�,  j   ��}j  �   U�  �   ��}�  �   ��}�  ]   ��}]  �   U�  ~   ��}~  �   V�  �   ��}�  �   U�  3   ��}3  5   P5  �   ��}�  �   U�  �   ��}�  �   U�  '   ��}'  >   U>  �   ��}�  �   U        ;  j   R�  �   R�  �   V�  �   p� ��  �   R�  �   V�  "   p ���"  4   R4  n   V�  �   R�  �   V�  �   r� ��      R      V     w���  +   R+  B   VI  T   RT  ]   V]  s   Rs  v   p ���v  �   p}����  �   w����  �   R�  �   V�  �   r��  �   w����  �   R�  �   V�     w���  D   RD  O   VX  f   R�  �   R   :   R:  A   VA  S   p ����  �   R�  �   p ����  �   ��}2����  �   R�  �   p ����  �   w����      V      p ���     v~���     ��}2���     V  '   p ���'  7   R7  ;   p ���;  b   r~���b  o   Ro  >   w���>  B   p ���B  J   ��}2���T  [   p ���[  `   ��}2���`  g   p ���g  l   ��}2���l  p   p ���p  �   ��}2����  �   r~���        g  �   V�  �   V      V$  0   V4  @   VD  P   Vh  �   VB  I   V     V0  9   VO  X   V     V�  �   V�  �   ��}�  �   V�  �   V�  �   ��}'  f   Vf  j   ��}j  o   Vr  y   V{  �   V�  �   V�  �   V�  �   V�  �   V�  �   V�  �   P�  �   V�  �   V�  �   P�  �   V�  �   V�  �   R�  �   P�  �   V  	   P	     V     P     V'  )   P)  .   V7  9   P9  >   V�  �   V        W  �   U�  �   V        �  �   V        �  �   W        �  �   P        �  �   �         �  �   R        �  �   V        �  "   ��  :  �   ��  �  �   ��  �  '   ��  >  �   ��          �  "   p�:  S   p�S  �   ��}�  �   p��  �   ��}�     p�     V     ��}  '   p�>  B   p�B  T   ��}T  [   p�[  `   ��}`  g   p�g  l   ��}l  p   p�p  �   ��}        �     W     R  "   W:  y   Wy  �   R�  �   W�      W      R  '   W>  �   W        �  "   � :  �   � �  �   � �  '   � >  �   �         �  �   �         :  M   �           '   �         �  "   ��  M  �   ��  �  �   ��        ��  >  �   ��          �  "   p�M  S   p�S  �   P�  �   p��  �   P      p�     V     ��}     P>  B   p�B  K   ��}K  T   PT  [   p�[  `   P`  g   p�g  l   Pl  p   p�p  �   ��}        �  "   ��}M  �   ��}�  �   ��}      ��}>  �   ��}        �     W     R  "   WM  y   Wy  �   R�  �   W      R>  �   W        �  "   p�M  S   p�S  �   ��}�  �   p��  �   ��}      p�     V     ��}>  B   p�B  T   ��}T  [   p�[  `   ��}`  g   p�g  l   ��}l  p   p�p  �   ��}        P  �   V�  �   V     VO  T   VX  `   Vd  l   V        
     P     p|�        �  �   P        �  �   Q�  �   qy��  �   Q        �  �   U        �  �   V        4  C   w�C  �   W        4  Q   QQ  S   qy�S  �   Q        G  g   Rg  �   w        4  �   U        W  �   U        W  �   �         v  �   P        }  �   V        �  �   R        �  �   �         �  �   Q        �  �   V�  �   r 2$� "             Q        ~  �   W        �  �   Qo  >   Q        �  �   Vo  r   Vr  y   u 2$� "
 y  {   V{  �   u 2$� "
 �  �   V�  �   u 2$� "
 �  �   V�  �   u 2$� "
 �  �   V�  �   u 2$� "
 �  �   V�  �   u 2$� "
 �  �   V�  �   u 2$� "
 �  �   V�  �   u 2$� "
 �  �   V�  �   u 2$� "
 �  �   V�  �   u 2$� "
 �  �   V�  �   u 2$� "
 �  �   V�  �   u 2$� "
 �  �   V�  �   u 2$� "
 �     V     u 2$� "
      V     u 2$� "
   '   V'  .   u 2$� "
 .  7   V7  >   u 2$� "
         �     U        �     r 2$� "
      q 2$� "
         �  �   ��}        f  �   P        f  �   Q�  �   qy��  �   Q        w  �   W        f  �   V        �  �   w��  �   W        �  �   Q�  �   qy��  �   Q        �  �   R�  �   w        �  �   V        �  �   V        �      �         �      Q        �  �   R�  �   v 2$� "        �  �   P        �  �   Q�  �   qy��  �   Q        �  �   W        �  �   V        '  4   ��}        4  b   ��}�  �   ��}        U  b   ��}        �     P  �   ��~�  �   �P��  �   P�  �   ��~�  �   �P��  =   ��~=  R   �P�R  u   ��~        �  ]   R]  �   ��~�  �   �R��  �   R�  �   �R��     R  =   ��~=  R   �R�R  u   R        �  �   P�  �   ��~     R!  &   R        �  �   0��  �   ��~�     ��~3  @   P@  �   ��~�  �   ��~=  R   ��~        �  �   ��~�  �   ��~��  �   ��~�  �   ��~��  =   ��~=  R   ��~�R  u   ��~          �   0��  R   0�          �   4��  R   4�          �   ��~�  =   ��~        ]  y   ��~#�y  �   P        y  �   W        ]  �   �2�          ]  �   P        ]  q   Qq  s   qy�s  �   Q        g  �   V        ]  �   W        �  �   ��~�R  l   ��~�l  u   P        �  �   PR  l   Pl  u   ��~#H        �  �   ��~R  u   ��~        �  �    [���R  u    [���        ^  l   ��~�l  u   P          "   P             ��~  "   W             ��~        <  c   �P�=  R   �P�        <  X   ��~#����=  G   ��~#����        r  v   Pv  �   v �  �   P        �  �   U        r  �   �p�          r  �   P        r  v   0�v  �   Q�  �   qy��  �   Q        �  �   W        r  v   0�v  �   U        �  �   P        �  �   ��~        �  �   ��~        �  �   P�  �   v �     P        �  4   U          4   P        �  4   �/�          �     P        �  �   0��  �   Q�  �   qy��     Q        �  %   W        �  �   0��  4   U          4   ��~          4   ��~        T  c   P        T  c   ��~        T  c   Q        L  T   PT  c   v         L  c   ��~�        z  �   P        z  �   ��~        z  �   W�  �   ��~        �  �   P�  �   v         �  �   ��~�        �  �   r ��        �  �   P�  �   v 2$� "�        �     P  &   ��~#�&  =   P        �  =   ��~          =   Q             R    
 p 2$� "�  &   ��~#�2$� "�&  ;   R;  =  
 p 2$� "�        �  �   P�  �   V�  �   �P�        �  �   R�  �   U�  �   �R�        �  �   �         �  �   �|        �  �   P�  �   P        �  �   ��~�p  �   ��~��  �   P�  �   p�  �   ��~�        �  �   Up  �   U�  �   �R�        �  �   Vp  �   V�  �   �P�        �  �    [���        x  �   ��~��  �   P�  �   p�  �   ��~�        x  �   V�  �   �P�        �  �   P�  ,   V,  .   �P�.  9   V9  ;   �P�;  D   V        �  �   R�  -   W-  .   �R�.  :   W:  ;   �R�;  D   W        �     P  .   P;  D   P        �  ,   V,  .   �P�;  D   V             Q  .   Q;  D   Q             R  '   R'  ,   p 2$v ",  .   p 2$�P";  B   RB  D   p 2$v "        P  o   Po  �   W�  �   �P��  �   W�      �P�      W        P  o   Ro  �   V�  �   �R��  �   V�      �R�      V        o  w   P�  �   P�  �   P�  �   P        o  �   R�  �   ��~�  �   R�      ��~        o  �   V�  �   V�  �   �R��  �   V�      �R�      V              P   �   V�  �   �P��  �   V�  �   �P��  �   V          1   R1  �   W�  �   �R��  �   W�  �   �R��  �   W        (  +   P+  1   v1  �   ��~        /  1   P1  �   ��~        1  V   P~  �   P�  �   P�  �   ��~�  �   R�  �   P�  �   P�  �   R        X  j   P�  �   P        1  �   :��  �   :��  �   J��  �   :�        �  �   U        �  �   W                 P    k    Uk   �    P�   !   U!  !   �P�!  m!   Um!  n!   �P�n!  �!   U�!  �!   �P��!  �!   U            &    R&   k    �R�k   �    R�   �!   �R�            &    0�&   f    P�   �    P!  U!   P�!  �!   P        A   R    WR   f    p 2$u "�   �    p 2$u "!  !   p 2$u "!  !   �D!  (!   p 2$u "        D   f    V�   �    V!  H!   V�!  �!   V        !  !   V        �   �    �\��   �    P        �   �    P�   �    r�         �   �    R        �   �     [���        �   �    �\��   �    P        �   �    4�        �   �    R        �   !   4�U!  �!   4�        �   !   U!  !   �P�U!  m!   Um!  n!   �P�n!  �!   U�!  �!   �P�        �!  �!   P        n!  �!   4�        n!  �!   R        y!  �!   Q        |!  �!   P�!  �!   r        �!  �!   ��!  �!   R�!  �!   ��!  "   R        �!  �!   V�!  �!   V�!  "   V        �!  �!   P�!  "   P"  "   r 2$q "         "  3"   �3"  P"   PP"  W"   �W"  s"   Ps"  �"   �        H"  R"   QW"  k"   Qk"  n"   p ["���s"  �"   Q�"  �"   [�"���        P"  R"   Ps"  �"   P        #  #   P!#  2#   P        �#  ,$   Q        P$  g$   � g$  |$   r |$   %   u %  �%   �         �$  �$   P�$  �$   P�$  �$   P%  %   P %  #%   Pd%  u%   P        B%  �%   ��|�%  �%   ��}�        �%  �%   P�%  �%   V        �%  �%   W�%  �%   q         �%  �%   � �%  �%   r �%  &&   u&&  f&   �         �%  �%   ��%  �%   r�%  &&   u&&  f&   �        �%  �%   ��%  �%   r�%  &&   u&&  f&   �        &  -&   P        9&  9&   P9&  ]&   V        9&  `&   W`&  f&   q         p&  �&   � �&  �&   r �&  !'   u!'  $'   �         �&  �&   P�&  �&   P        �&  �&   P�&  '   V        �&  '   W'  $'   q         0'  _'   � _'  t'   r t'  �'   u�'   (   �         �'  �'   P�'  �'   P        �'  �'   P�'  �'   V        �'  �'   W�'   (   q          (  .(   � .(  =(   r =(  �(   u�(  �(   �          (  .(   �.(  =(   r=(  �(   u�(  �(   �        O(  Y(   PY(  s(   W�(  �(   P�(  �(   W�(  �(   W                P   A    P            	    R	   @    U@   A    �R�            	    0�	   !    Q!   #    qy�#   A    Q           /    R/   =    p            	    0�	   ?    W?   @    u @   A    �R        p   �    P�   �    t �   �    �`�   �    t �   	   �`	  #   t #  '   �`'  ;   t         p   ~    R~   ;   �d        ~   �    R�   �    V�      R     �l'  ;   �l        �   �    W�   �    V�      W'  ;   V        �   �    P        @  N   PN  �   �h        @  d   Rd  �   �l        X  �   U�  �   � #�        X  �   V�  �   v�        _  x   Wx  y   t y  �   �P�  �   w��  �   W�  �   V�  �   v��  �   V        �  �   P        �     P     �P�  ,   P,  5   �P�5  H   PH  J   �P�J  U   PU  W   �P�        `  v   Pv  �   �P�        `  �   R�  �   �R��  �   R        �  �   P�  �   �P��  �   P�  �   �P�        �     R  G   �LG  V   RV  [   �L[  g   Rg  l   �Ll  x   Rx  �   �L�  �   R�  �   �L�  �   R�  �   �L�  �   R�  �   �L�  �   R�  �   �L        �     �   D   VD  G   PG  Y   � Y  [   V[  j   � j  l   Vl  �   � �  �   P�  �   � �  �   V�  �   � �  �   V�  �   P          G   RV  [   Rg  l   R�  �   R�  �   R�  �   R        �  �   V        �  �   Q�  �   qy��  �   Q        �  �   R�  �   v        �  �   U        �  �   � �  �   V�  �   v|��  �   p|�        #  '   P'  y   W        �  �   P�  �   V�  �   �P��     V     wv�  Z   �P�Z  �   V        �  �   W�     W     w�  4   W4  E   w�E  Y   WZ  �   W        �  �   Q�  �   Q�  �   P�  �   R�  1   R1  <   q�?  B   PB  Z   RZ  �   Q�  �   P�  �   R        �  �   Q        �  �   q        �  �   R        �  �   r        �  Z   �)          �     R        �     r        �  �   P�  �   U�  �   �P��  �   U�  �   �P��  �   P        �  �   R�  �   V�  �   V�  �   V        �  �   0��  �   Q�  �   W�  �   Q�  �   W�  �   Q�  �   W�  �   0�        �  �   0��  9   �\�  �   �\�  �   �\�  �   �\�  �   �\�  �   0�        �  �   0��  �   �P�     P  �   �P�  �   �P�  �   �P�  �   P�  �   �P�  �   0�        �  �   0��     �T     P  �   �T�  �   �T�  �   �T�  �   0�        �  �   W�  �   Q�  �   W        Z  x   Px  �   R        �  �   V�  �   V        �  �   V              P  &   U&  '   �P�              R  '   �T           *   � *  $   V           C   0�C  �   �L�  �   Q�     �L          �   W�  �   P�  %   W        *  .   P.  '   �P        �  �   Q�  �   �L        �  �   P�     R        C  W   v        ]  n   �T        ]  n   V        �  �   V        n  t   V     V        �	  �	   P        �	  �	   P        �	  �	   W�	  

   �        �	  �	   V�	  

   �        �  �   � �  �   p        �  �   ��  �   P        �  �   ��  �   p        �  �   ��  �   Q        �  �   ��  �   Q        �  �   ��  �   p        �  �   ��  �   P        �  �   � �  �   p        �     �   7   p        �     �  7   P        �     �  7   P        �     �   7   p              �  7   P              �   7   p        d  �   P        d  �   V        d  �   0�        �  �   � �  �   R�  �   p        �  �   ��  �   P        �  �   ��  �   p        �  �   ��  �   p           $   � $  -   R-  K   p           $   �$  K   P          $   �$  K   P        f  {   � {  �   R�  �   p        �  1   � 7  �   �         �  �   @[��  �   r��     <[�  ,   R7  C   r�C  E   Rh  �   R�  �   @[�        �  ,   0�,  7   P7  h   0�h  �   P�  �   �l�  �   0��  �   P        �  �   P�  �   �           �   V�  �   U�     U     V        �  <   0�<  A   PA  �   U�  �   P�  �   0��     P        U  \   p ��\  a   Pa  h  
 v�3%��i  p   P        ^  i   U        �  �   <[��  �   <[��  �   R�  �   <[��     R        ���        ������Ց����        p�s�w��        ��В���        �������        +�/�3�������        @�������        ����#�� ��        G�S�V�j�        ����Д�        "�'�,�1�9�K�`����        `�f�k�q�        ��G� ��/�I�K�Q�        ����ĖƖ        ��ĖƖ���        ������        ���7�        N�R�[�u�Й���        V������        �0�0�{�������� �������� �� ��        ��        $�)�-�6�e�p�        6�M�Q�`�         �p�p�ӛ��6�        @���        ؜ۜ��        h�{�����        m�{�����        m�p�t�w�        ��ȞО�����f�        Ҟ՞ڞ���        ���>�C�H�X�        ����        !�$�)�3�C�H�        ~�����ݟ�^�        ��ȟ˟Ο        ��6�;�@�P�        �������        ���(�;�@�        l�y���Y�        ��������        ǠʠϠ�        ��1�6�;�K�        ������        ���#�6�;�        r����I�        ��������        ������֡        ֡��!�&�+�;�        �����        ��	��&�+�        `�k�p�u�        ãƣˣۣ        �����������ˤD�        �!�&�3�        ˤФ��1�6�        ������        ���#�6�=�        ;�>�C�P�        P�������        ��������        V�Y�b���Х� ���        r��� �j����        r��� ��        ~��� ��        ���
�        � �%�E�        E�j����        P�S�V�e�        ������������        ����Х�        ӥ֥ۥ�        ƦɦҦJ�`�{����        ��	��        ����էߧ        ��������        ������ǧ����        �J�`�{�        c�f�k�{�        +�@�`���        2�6�����        6�@�`���        J�N�S�`�        ި� �� �J�        ި� ���� �J�         �� �J�        ��E�J�        �� �E�        y�}����        y�}����        ����        ��
��        &�)�/���Ӫ���� �        ?���Ӫp�����        U���#�p�����        <�?�D�T�        u����� �P�v�{�����        u�֫��� �P�v�{�����        u������ �P�v�{�����        ��ά �P�v�{�����        ��������v�{�        ��ά �P�����         �P�����        ������֫        ������ѫ        ����īѫ        ������ī        �p�� �P�v�{���        �F�� �P�v�{���        ��� �P�v�{���        ��P�v�{���        ����q�v�        ���P�q�{���        P�q�{���        ���-�F�        ���-�A�        ���2�A�        ��-�2�        H�K�P�p�        Ӫ���        ���#�        ��ŭ���        ������ŭ        Эӭح���        ����p���        s�v�{���        ������ʮ        ���*�        ���*�        M�h�p���        r�u�z���        ������[�p�˰���        ��*�p����\�t���        ���p����7�        ̯ԯ"�)�        ԯ�p����"�)�7�        p����"�)�7�        s�u�x�~�)�7�        ~����"�        ���*�        7�\�t�y�        B�E�H�W�        ������������        *�[���˰        ������˰        ���˲�;�P��        /���� �P�̳��        /���� �P���        <�D�����        D�Z�� �P�������        � �P�������        ��������        � �P���        ��������        ��̳��        ������ǳ        ���������        ��˲ �;�        #�&�+�;�        b� �0�����n�        u��0�p����4�n�        u�մ0�p�����        ������        ����0�p�������        0�P�������        3�5�8�>����        >�P����        ������ϴ        ״ڴߴ�        ���4�9�        ����        D�G�L�V�`�g�        � �p���        s�v�{���        ������G�`���з��        ���`���зL�d���        ����`���з'�        ������        ��ֶ`���з��'�        `���з��'�        c�e�h�n��'�        n���з�        �����        '�L�d�i�        2�5�8�G�        t�w�|�������        �G�����        ��������        Ÿɸ̸w���� �κ        ۸F���й �|���κ        ۸,���й �W�        ��B�I�        ����й �B�I�W�        ���� �B�I�W�        ��������I�W�        ���� �B�        .�1�6�F�        W�|�����        b�e�h�w�        ����������Ǻ        F�w�й�        ӹֹ۹�        ������������ ��        �p���� ������        �V���� �w�        ��b�i�        �0���� �b�i�w�        ��л �b�i�w�        ��������i�w�        ��л �b�        X�[�`�p�        w�������        ��������        ļǼ̼ּ��        p�����        ������        &�)�/���K�`�.�        ?����0�`�ܾ��.�        ?����0�`���        L�T�����        T�j��0�`�������        ��`�������        �����������        ���`���        ��������        ��ܾ����        ¾žȾ׾        ���� �'�        ���0�K�        3�6�;�K�        F�I�O����k���N�        _�ʿ�P������N�        _����P�����        l�t�����        t����P���������        �0���������        ��������        �0�����        ������ʿ        ������        ��������        $�'�,�6�@�G�        ʿ��P�k�        S�V�[�k�        ����������ϜМ�� ���5�@�ƝН���� �� �;�@�����f�p�^�`�Y�`�I�P�u�����u�����D�P�������� ���������ŨШJ�P�e�p�����ש�� �� � � �?�@�_�`����Ү�2�@������������� � ���� �%�0�>�@�E�P�n�p�~�����������κкպ����� �� �.�0�5�@�N�P�U�        ���#�/�        B�G�Z���        ������        +�;�>�P�        0�;�>�P�        P�`�c�h�        }�������        ��������        +�@�`���        2�6�����        6�@�`���        ����`�v���������������/�0�@�@���������� �i�p��� �� ������� ��        ��"�~��������        ?��������������        S�b�_���        b�p������_���������        b�p���� �@�����        b�p���������        ��������        ���������� �        ���������� �@�        ����������        ��������        ���@�W�����        ���@�O�        ������        ������������        ��������        ��������        ��$�2����        ��������        ��������        i�l�q�~�        )�U�`������        d�U�`������        d�R�`�����C�f���        ���f�z�        ������������C�        �����������        ����������������        ������
��        �����������        �������������C�        ���������.�        ��������        ��z���        R�U�I�L�Q�f�        �������        ��������        ����������        &�)�,�0�@��        D�������@�Y�p������        J�M�a�i�l�q�        ��������|���        ��������        �����������p�P���P���|�        '�*�-�t�p����P���0�        p����P���0�        ���������P���0�        �������������P���0�        �������������P���0�        ������������        ����������������0�D�        ����������������        )�B�D�X�[�t�        )�7�D�S�        7�B�e�t�        ��������P���P���        R���P���        R�`�l���P���        R�`�w���P���        ��������C�F�N�Y�        ���������        ��������        &�)�,�p�{�x�        {�� �M�Q�a�p��������        {�������        {�~�����        ������������        ��������������        ��������        �� �-������� �5��p���`�����        �� ������5�L�`�        �� ���L�[�        �� ���        �� ���        �����5�        �����&�        Q�T�W��� ����p���L�         ����p���L�        0�3�:���0�p���L�        0�3�B�������0�p���L�        0�3�M�������0�p���L�        ������������        ��������        �������        �������         ���"�p��p���        r��p���        r������p���        r������p���        ���������������Q�T�V�a�        �����-�        ��������        <�?�D�N�c�j�        ������������        �������������������        ����� �(�����L�����        ����������#�L�����        ����-�L�        ����-�@�        #�-�����        ��� �E���        ��� �E�W�\�_�        q�t�y�{�~���        {�~�����        �� �����        � �����        �����������        ��������        ������        ��������        ���0�        R�U�Z�d�{���        ��������        �� �� �� �x�����        ����        ��������        ������f�p�������        ��������        �������        �L�p�z���������        +�.�0�8�        L�Y�����        L�R�����        R�Y�����        Y�f�����        Y�_�����        _�f�����        8�P�V�n�        x�������        �������        ��%�9�E�M�_���        ��+�5�        ������ �        ��������        )�9�E�M�        )�,�/�2�        ,�/�2�9�E�M�        ������� �{�        P�S�W���������H�        P�S�W�����H�        P�S�W�`�m�����H�        Q�S�W�Z�]�_�l�o�r�u�        ��������������������        ����������������        ����������������        A�C�G�J�M�O�U�X�[�^�        ��������������������        ����������������         �$�(�,�9�<�G�J�        ����������������k�|�        ����������������        ����������������;�L�        ����������������        P�T�X�\�b�h�        ����������        ��������������������        ��������������������        1�3�7�:�=�?�L�O�R�U�         ������'�*�        a�c�k�n�q��������)�        a�c�k�n�q�s�����        0�4�8�<�B�H�        ������������        ����������������        ������%�+�        q�s�{�~���������        ������ �        ��������        PTX\bh        ������        ������        @DHLRX        bdgkoqw}        ��������        ��������        ��������        ACKNQdgj��        ACKNQSY_        �.	2	<	        ]	�
�
�        �	�	�	`
�
�
 d��        �	�	�	�	 S��        �	�	�	
�
�
��        �	�	�	�	  d�        �
�
�
 ��        �
 ��        	$��        P`=?AZ $        FU $        `�w�@p��
        `q}��@Ucp
        `q��@U
        ��@I        }cp        q}�w�Uc��        w���        �=?A� $@���
        �������
        ������        �� $@        =?A        7��x        ���x        ����� Jx        ��� `x        � `i        ��J`        ���� J                 ����        �        #^bl        |��0�        ���0�����        ����        ����        ��������        ����        ������        ����        ���         #2P�         #&        &2P�        PVX[        U~�        ����0@        ����0@        ����        ����@P        ����        ��@P        �'Pp        -58>         058>         S|0P        ���� 0        ����        �� 0        ����        ��p�        ���J����        JMV��        ��        NR\        c���        �Q`��7         ��         ���         ��        Q`����#^s�7         A��        GORXp�        JORXp�        m���        ������        ����        ����        ���        
                  0Y`�        gjm{ 0        gjmp        p{ 0        ��@`        ����P`        ����P`        �� @        !`p                !`p        'S          Yadj0@        \adj0@        ��         ����@P        ����        ��@P        ����        ����         Q`}��        C ~ � �         � 1$@$k$�$(        � � �%�%        � � �%�%        � � �%�%        � 1$@$k$�$�%�%&�&'>'S'�'(        � !!�%�%        '!/!2!8!P&`&        *!/!2!8!P&`&        M!v!�%�%        �!�!�!�!`&&        �!�!�!�!        �!�!`&&        �!�!`%�%        �!�!�!�!�% &        �!�!�!�!�% &        "9"@%`%        G"J"M"[" &&        G"J"M"P"        P"[" &&        a"�" %@%        �"�"�"�"0&@&        �"�"�"�"0&@&        �"�" % %        �"�"�"#@&P&        �"�"�"�"        �"#@&P&        #3#�$ %        9#A#D#J#& &        <#A#D#J#& &        _#�#�$�$        �#�#�#�# &0&        �#�#�#�#        �#�# &0&        �#�#�$�$        �#�#�$�$        �#�# $1$@$]$`$k$        #(^(b(l(        s(�(�(�(        �(�())        4)-*@*�*        T)[)])g)`*�*        �)�)�)�)�)�)        �)�)�)-*        �)�)�)*        �*�*�*�*        +>+B+L+        S+�+�+�+        �/�/�/.1@1S1        �0�0�0�0        1�1�1�1        �1�1�1�1        e2�5�5^:        e2k2l2o2        t2{2~2�2�8�9*:^:        �8�9*:^:        �2�2�23�5�5�5�6�7�8         6�6�7�8         6#6'6�6�7808�8         6#6'60686�6�7808�8         6#6'606C6�6�7808�8        3�5�6�7�8�8�9*:        `3
4�9�9        b3e3g3{3}3�3        �3�3�3�3        �3�3�3�3        �3
4�9�9        �3�3�9�9        4(4+4.4        K4N4T4W4Z4b4e4h4        �4�4�4�4�6P7�9�9        �4�4�4�4�6P7�9�9        #5+505A5        A5f5�9�9        f5t5�9�9        i5t5�9�9        �5�5�5�5        �:�=�=~B        �:�:�:�:        �:�:�:�: A�AJB~B         A�AJB~B        �:�:�:6;>>>�>�?�@         >�>�?�@        @>C>G>�>�?0@P@�@        @>C>G>P>X>�>�?0@P@�@        @>C>G>P>c>�>�?0@P@�@        >;�=�>�?�@ A�AJB        �;*<BB        �;�;�;�;�;�;        �;�;�;�;        �;�;�;	<        <*<BB        <<BB        4<H<K<N<        k<n<t<w<z<�<�<�<        �<�<�<
=�>p?�A�A        �<�<�< =�>p?�A�A        C=K=P=a=        a=�=�AB        �=�=�A�A        �=�=�A�A        �=�=�=�=        �B�B�B�C�CTD        �B�B�B�B        �B�B�BC        �B�B�BC        CNC�C�C�C�C�C D        qCtCwC�C D.D        qCtCwCzC        zC�C D.D         DDDD        �D�DEGENE�E�EG        EEEE        `E�E�E�E FG        lEsEuE{E FIF�FG         FIF�FG        �E�E�F�F        !E,E.E3E        7E;E?EGENE`E        �E�E�E�E        �E�E�E F        TGYGeG�G�G�G        �G�G�G�G        �G�G�G�G        HH HNI`IK        HH HCH@JMJPJ^JaJ�J�JK        @JMJPJ^JaJ�J�JK        QJ^JaJ�J        VHXH[H^HaHdH        MJPJ^JaJ        /K|KK�K�KsLvLyL�L�M        /K2K4K7K        9KaKdKgK        �KsLvLyL�L�M        �K�K0M=M@M�M�M�M        0M=M@M�M�M�M        �KsLvLyL�L0M�M�M        �K�K�K�K�K�K        �KLLL         LBL�M�M        �L�L�L�L        �N�N�N�O�OXQ        �N�N�N O�P�P�PQ$QXQ        �P�P�PQ$QXQ        O O#O&O        �O.P2P:P        �R�R�R SSS
S�S        SSS]S        SSS#S        �S�S�SU0U�V        �S�S�S�SVV V.V1V�V�V�V        VV V.V1V�V�V�V        !V.V1VkV        TTTT        PU�U�U�U        V V.V1V        �W�W�W�X�XHZ        �W�W�W�W�Y�Y�Y�Y�Y�YZHZ        �Y�Y�Y�Y�Y�YZHZ        �Y�Y�Y�Y        �W�W�WX        �Y�Y�Y�Y        [)[@[�[�[(\        @[�[�[(\        <\Y\p\]!]X]        p\]!]X]        l]�]�]^^S^        �]^^S^        f^k^�^�^�^�^�^` `;a        +_f_�`�`�` a a;a        X`�` a a        �a�a�a�a�a/c@c[d        Eb�b�cdd d@d[d        xc�c d@d        �d�d�d�d�d�d�de        �d�d�d�d        e/eSese�e�e�e�e        Se[e�e�e        /eAese�e�e�e�e�e        se{e�e�e        	fafcfffpfi        )f,f0f7f:f@f         g�g�h�h        gggggg        gggggGg        Gggg�h�h        Qg`g�h�h        �g�g�h�h        �g�g�g�g�g�g�h�h        �g�g�h�h        h�h�hi        ,h/h;hDhFhHh        �h�h�h�h        iii�j�j�jkm        iiAiDiIiSi        �k�k�k�k�k�k        �k�k�k�k�k>l        �i�i�j�jkDk�k�k        �i�i�i�i�j�j�j�jk3k:kDk        �i�i�j�j�j�jk3k        �j�jk k        �i�i:kDk        �i�i�i�i�j�j�j�j3k:k�k�k        �j�j�k�k        �iOj�j�jkk�k�k�l�l        �i�ikk�k�k�l�l        kk�k�k        �iCj�j�j        �i�i�i5j7jAj�j�j        OjojDkXk        YjhjDkXk        ClFlLlfl        �l�l�l�l        mm)m�n�n(o        mm)m,m        |m�m�m�m        Onnn�n(o        On\n`nbn�n�n�n(o        On\n�n�no(o        �n�noo        `nbn�no        \n`nbnnn�n�n        �n�n�n�n        :oAoOoJq`q�q        :oAoOoRo        �o~p�p�p        q7qsq�q        q%q)q+qsq�q�q�q        q%qsq�q�q�q        sq�q�q�q        )q+q�q�q        %q)q+q7q�q�q        �q�q�q�q        r�s�s�s�s=        #r+r-r<r        Pr�r sust t�}$~        Prcrnrpr s=sRsWst t        Prcr s=st t         s)stt        nrprRsWs        crnrpr�r=sRsWsus�}$~        `sls�}�}        �r�r tPtdu�u        �r sPt�t�tuPudu�u�}$~�~�~         �r�r�r�r�t�tPudu$~<~        �tu�u�}<~�~�~         v&v�~�~�~�~        �y@{�~         GzXz�~        rz�z         Pvfv^~�~�~�~        �x�x }�}        <y@y�}�}        ^tftht�t�~�~        �s�s�s�s�t�tu6u&*        �t�tuu        �t�t�~�~0=        �t�t�~�~        W��^�        �����^�        ��������6�^�        ������C�^�        ��C�L�        ��6�C�        �����6�        ����        w���~�        ������Հ�~�        ������ƀʀ̀��V�~�        ������ƀ��c�~�        ��c�l�        ʀ̀V�c�        ƀʀ̀Հ�V�        ��'�0�        ������Ԏ�'�        +�6���S���������W���        +�����6���S���������W���        ^�f�؆� �@�        ^�f�0�@�        ^�f�8���������@�        @���������@�        f��������C�@���        f�z���������������p���        f�z���������p���        ����p�|�        ������        z������������������C�@�p�        $�0�@�L�        Ђ��0�l���        �����������C�]� �`�        �����������Ѓ݃�C�O�R�U� �0�        ���������ЃC�O�R�U� �0�        C�O� ��        ��݃�        �����Ѓ݃����O�R�U�]�0�`�        ���0�<�        ���]� �����`���=�F�        �5�]���`���        ����`�l�        [�������        ��������        �����������        �������        ���0�0�        ��׊0�t����� �0�        ��Ɋˊ0�H�U�Z�����        ��0�H�����        0�<�����        ɊˊU�Z�        Ɋˊ׊H�U�Z�t� �0�        c�o� ��        �������        ��̋�� �        ��ŋ�� �        ��؆0�V�.�=�        Ɔ҆0�<�        ���� ��.�        ���.�        ،܌}���        F�R�U�X�        W�c�f�i�        \�_�b�p���        \�_�b�e�        e�p���        p���̎Ԏ        v���̎Ԏ        ��W�����        ������        ���"�        '�C�I�W�        1�<�I�W�        ��ЅӅօ        ����        )�,�/�9�<�?�        9�1�@�����ל        ۏ�@��C�C�N�i��X�        ۏK�g��@��C�C�N�i��X�        ������Е�        �����        ���0�3�6�P��        �0�3�6�P��        �C�C�`�����P�        �*�5�7�C�O�R�U�Ɣ˔ �P�        �*�C�O�R�U� �P�        C�O� �,�        5�7�Ɣ˔        *�5�7�C�O�R�U�`���Ɣ˔�� �        Ԕ�����        ����͘���C�        ����e�g�n�����đ�����        ��������e�g�n����������������        ����e�g�n������������        �������        ��������        ������������������đ��������        �������        ɐL��ЕP�p��;����        ɐ��P��;�        3�?���        �I�P�p�        >�I�P�p�        L�e�g�n�p���        V�e�p���        P�͘����        `�����$�C�`�����        `�r�y�{������
�C�`�        `�r�����C�`�        ���C�K�        y�{��
�        r�y�{������
�$�����        ������        ��������        `�|�����        j�u�����        `������ޚ�        v������        ��������͚ޚ        ����͚ޚ        ����-�O�        �����        ����        ��� �����        ����        � �����         �1�|���        &�1�|���        i��X�c�        ��������        ��ɛϛқ        כ����        �����        f�������        ������        ٓܓߓ���        ������Z�p�̝        D�G�L�Z�����        D�G�R�Z�����        ��������        ٝܝߝS�`�v�        ٝܝߝ�        )�,�/�2�        <�?�B�H�M�S��@�        B�H�M�S��@�        ����        ��������        ������Ğ        ��������        ʞ�@�A�F�X�        ������̠��+�u�        ��������         �@� ���K�W�         ����        �"�(�1�        ��П������Ĩ�0�<�?�F�������        ��П��������������Ĩ������        ��������        �������������0�<�?�F���        ��������<�?�F���        ����M�i�        ����M�`�        �����0�        ҟٟզ�         �y�� �0�`�������        �����        ���5�0�F�        �(�/�5�0�?�        �(�/�5�        %�(�/�5�        5�Y��0��� �F�`���        5�A�D�G�K�M���ܢ� �F�`�        5�A�D�G���ܢF�`�        5�A���̢        K�M�� �        A�D�G�K�M�Y��0�ܢ���        �����        a�~��������� ��        a�p�s�u�        ��������        "�I���������`�v�        0�<�C�I�`�o�        0�<�C�I�        9�<�C�I�        I�q����v�������        I�U�X�[�c�e���ơv���        I�U�X�[�v���        I�U�����        I�U�����        c�e���ơ        U�X�[�c�e�q�����ơ�����        ϡۡ����        2�o�ФХ��Ӧ���        Q�T�W�c�g�j�        ��� �        �� �=�Щ�        '�6�Щ�        X�z���ĥ��¦        X�g�j�l�        ������ĥ        ����        +�.�0�2�        o�����$�0�Х�        }�������Хߥ        }�������        ��������        ����0�p��0�`���        ������������A�E��0�        ���������0�        ������        ����� �        ����A�E�        ������������0�A�E�p�`���        N�Z�`�l�        y�|�������        y�|�������        y�|�������        ������̠��        ��̠��        f�i�m����� ���0�<�?�F�        x�������0�<�        x�������        ��������        ��� ��        ������2�C��        �
�C�����ͫ        ��� ��C�P�`�z�~���        ���C�P�`�z�        C�K�`�n�         ��~���        �� ��
�P�`�z�~���ͫ        P�X�����        !�$�'�2�����        !�$�'�*�        *�2�����        ��������        ����������[�        X�z��� � �=�        X�l�p�r�����Ь�� �        X�l�����Ь�        ����Ьެ        p�r�� �        l�p�r�z���Ь�� �=�        ��Ȭ �,�        �������� � �        ��������        ���� � �         ����        f�i�l��#�ˮ        ȭ�#�p�����        ȭܭ��#�0�@�Z�^�p�        ȭܭ#�0�@�Z�        #�+�@�N�        ��^�p�        ܭ���0�@�Z�^�����        0�8�����        ����p���        ���
�        
��p���        p�v�x�{�        ܮ��#�0���        ������        �$�)�,�        2�>�D�G�        �A��������        ;�A��������        J�M�R�v�������        ]�i�p�v�����        ]�i�p�v�        f�i�p�v�        v����=���� �P�        v������������#����        v����������        v�����̲        v�������        �����#�        ��������������#�=� �P�        ,�8� �,�        P������        ����������`�v�        ��������`�o�        ��������        ��������        ��س��0�v���P���        ����óƳγг��v���        ����óƳv���        ����}���        ����}���        γг��        ��óƳγгس����0�P���        �"�P�\�        E���� �        _�k����        ���������#�        �������#�        �!�$�'�        *�J���        4�C���        ��̶Ӷٶ        u����ɻ        ̸ϸܸ�        ����ļ        ]�?���������0�h���        ]���������8���h���        ]�t��������8�[�g���        ]�t����8�[�        ���8�A�        ����g���        t��������������[�g�h���        ����h�q�        �����8�����        ������        ��������0�        ���0�        ܼ���3�@���        ������        �$�)�,�        2�>�D�G�        �8���ÿ`�p�        2�8���ÿ`�p�        B�E�J�n����p���        U�a�h�n�p��        U�a�h�n�        ^�a�h�n�        n�����$��������        n�z�}��������
�����        n�z�}�������        n�z�����        n�z�����        �����
�        z�}������������
�$����        ������        0�x�����        x�����������@�V�        ��������@�O�        ��������        ��������        �������V���`���        ����������������V���        ��������V���        ����]�|�        ����]�p�        ��������        �������������������`���        ���`�l�        ,�`��� �        F�R�����        �������+�3�        �����+�3�        �!�$�'�        :�Z� �+�        D�S� �+�        ��������        |���������.�        ��������        ��������        ��������        ����@�c��� �        ����@�c��� �        ����������� ��        �� ��� ��        �� ���        �� ���        �5������`�p���        ����'�)������`�        �����`�        ��!�<�        ��!�0�        '�)�����        ���'�)�5���������p���        ����p�|�        �� �c�h�         �#�`�c�h�l�����        
���#�����        
���#�        ���#�        #�G�l�����0����        #�/�2�5�=�?�}�����0�        #�/�2�5���0�        #�/����        #�/��� �        =�?�}���        /�2�5�=�?�G�l�}��������        ��������        ����`���        ����`�l�        ����������������        ������������        ��������        ��������        ��������        P�\�c�i�        ���0�3�@���        	����        4�D�I�L�        R�^�d�g�        ,�X�����p���        R�X�����p���        a�d�i���������        t�����������        t�������        }�������        �����<������� �        �������������"�����        ������������        ��������        ��������        �����"�        ��������������"�<��� �        +�7�����        @�������        ������������P�f�        ��������P�_�        ��������        ��������        ������ �f���`���        ���������������f���        ��������f���        ����m���        ����m���        �������        ����������������� �`���        ��`�l�        D�p����        ^�f�����        ������+�3�        ����+�3�        0�A�D�G�        :�Z� �+�        D�S� �+�        ��������        ��N�P�S�        ������i�v���        ��������        &�6�;�>�        D�P�V�X�        x�&��� �����        &�M��������� �6�        4�@�G�M� �/�        4�@�G�M�        =�@�G�M�        M�u�����6�������        M�Y�\�_�g�i�����6���        M�Y�\�_�6���        M�Y�A�\�        M�Y�A�P�        g�i�����        Y�\�_�g�i�u�������������        ��������        ����6�s�0�@�        ����6�@�        ����@�s�0�@�        ����������������@�V�        ��������@�O�        ��������        ��������        �����0�V����@�        ��������
�V���        �����V���        ���]�|�        ���]�p�        ���
�        ���������
�0��@�        ����        !�6�s�������        s������        ������������a�i�        ��������a�i�         ����        ����P�a�        ����P�a�        ��#�%�        �������������L�        ������������        ��������        �����        �������        ������        9�<�@�d�%�(�4�<�����        K�W�^�d�����        K�W�^�d�        T�W�^�d�        d���<�l��������        d�p�s�v�~���M�R����        d�p�s�v����        d�p�����        d�p�����        ~���M�R�        p�s�v�~�����<�M�R�l�����        [�g�����        @�S���p�s�w�        S�z�p�s�w�����        a�m�t�z�����        a�m�t�z�        j�m�t�z�        z�������P�0�`�        z����������������P�        z��������P�        z����,�        z���� �        ��������        �������������������0�`�        ����0�<�        t����@�        ������        ����������������        ������������        �!�$�'�        �,�����        �%�����        ��������        ����������������������������� �,�0�;�@�S�`�s��������������������������������� �!�0�?�@�O�P�_�`�o�p������������������������� �F�P�v�������������6�@�f�p���������=�@�����
��+�0�K�P�q�������������+�0�Q�`���������������1�@�a�p�����������+�0�?�@�a�p������ �;�@�O�P�q�����������0�0�n�p���������������� �H�P���������>�@�b�p������� �S�`������ �B�P���������<�@�����������2�@������� �S�`���������8�@������ �����|���L�P�i�p���������	��P�P���������)�0�{�����������3�@������� �S�`�)�0�I�P�����������H�P�������������&�0�j�p�������a�p�J�P�j�p�����������������' 0 w � ��LPip������� 8@x���� 8@Y`������� ,0;@GP]`��x������ $0;@��<	@	�  x��� lp��\`��7 @ � � ( (l(p(�(�())�*�*�* +L+P+�+�+�+�+9,@,�,�,�,�,)-0-y-�-�-�-. .i.p.�.�.	//Y/`/�/�/S1`1�1 252@2^:`:~B�BTD`D�D�DG GOGPG�G HKK�M N1N@N�N�NXQ`Q�Q�QRR�R�R�S�S�V�VW W�W�WHZPZ�Z�Z�Z [(\0\X]`]S^`^;a@awa�a[d`d�d�dee�e fiimm(o0o�q r=@^�`�~���'�0�ל��̝Нv���u�����[�`�ˮЮ����׷�\�`�ļм��������l�p�.�0�g�p�������������\�`���������� �����L�P����������        �� �"�0�2�@�B�P�R�`�b�        "�$�@��������� �        "�$�@�M�        ��������� �        "�$�@�������        "�$�@�M�        ��������p�������������� � � ���        ��:�G�[�        @�G�[�������        @�G�[���        ��������9�        �������        ��9���-�N�        ��9�>�J���        �������        ��������        ���o���        �*�6�v�        ���N�o�        ��������        ��������        �������        W�^�a�h�s���        i�e�s���        i���s���        i�r�t�z�        ��������        ��������        ����������O�P���        �������        ������������        <�G�P�������        C�G�����        P�_�����        "�%�0�N�        ��������        ����+�0���������i�p�� �*�0�:�        K�O�S�e�s������ �\�        Y�e�@�E�G�K�        s������ �@�        �������� �@�        ��������        ���� �)�        ��������        @�\�        ��������        ��'�0�8�@�G�        �'�0�8�        ��� �        0�3�5�8�        ��������        Y�\�b�m�����        Y�\�b�e�        e�m�����        ��������        �������        �����������        ��������        �������        ��������        ��)�H�K�Q�p���        ��0�;�p���        ��0�3�        3�;�p���        p�v�x�{�        ;�H�K�Q�        H�K�Q�_�        �������������0�        ���������0�        ��������        �����0�        ����        ��������        ��������        Y�������        Y�\�i�������        Y�\�p�{�����        Y�\�p�s�        s�{�����        ��������        ��@�P�p�        ����	�.�P�p�        ������P�p�        ������        ��P�p�        P�V�X�[�        ��������������         ����������         ��������        ������         ��������        ��������        ��������        I � � �         I L ` � � �         I L g r � �         I L g j         j r � �         � � � �         n��N        ����        ����        ������        �����         ����        ���         ����        ����        ����        ����                 ����        P`�                 ����        ����                ?�������        RX[^fi        ����        ���        ��        =@C�        =@CF        RXZ]                                $'),        ����        ����        ����        ����        ����        7:=AE��e	        7:EJY]        =AJW        ���e	        ����        ����        �	�	�	B
P
�
        �	�	�	�	        �	B
P
�
        �	
P
`
        

P
`
        �
�
�
�
        �
�
�
        �
�
�
        $        ���/2@        ���/        /2@F        ����        �����c��        �����        02        02        02        ORTW        ����        SV~���        VYfmp~����:        VYfmp~����        ����        ����        ����        ����        ����        ������        ����        ����        ����        U`�        &9<=        &6<=        9<=DGJ        DGJU��        DGJM        MU��        ����        `svw        `pvw        svw�        ����        ����*        ����        ����        ����                 ?BEY        BEf���        BEf�        ����        lo|���        lo|�        ����        /25I        KQ_{~���8        KQ_{~���        ����        ����        ����        ����        \_{~��        ����        �������n��        �������$        $';=        $';=        $';=        Z]_b        3Pp         Pp                 Pp        PVX[        ���n        ����        ����        ������        ����          ����        ��                   ����        ����        ���          #&<        uy}��        uy}        uy}        uy}        ����        � ��         $@Cw         $@Cc        [^r�        [^r�        /ps���        ���Cw        ����        ����        ����        ����        � CM        KNbil� 6        KNbil�        ����        ����        ����        ����         ����        ����0        ��0        ��0                N��.        fy|}        fv|}        y|}���        ������        ����        ����        ����        ����        ����        ����        ����        59=?Bj        59=?        59=?        59=?        X[]`        `���������G���ҀP���������������0�0�B�P���������p�p�����     2 @ � � � � �  Z`NP��� ����00� ;@ e	p	�
�
bp����kp��� ��00�  ``��ppx�np���� ��x�008@.0p        ���         Y ] c f i 6!@![!^!a!p!�!        �!�!�!�!�!�!        �!�!�!�!        @!F!I!L!        "4"<"]"        �"�"�"�"�"�"�"�"        p��  A P �! "f"p"�"�""#0#K#        `#�#�#�#�#�#        �#�#�#^$b$i$        �#�#�#�#        �#�#�#�#        �#�#�#�#        P#�#�#i$        �$�$�$U&p&�&�&9'        +%>%@%C%        >%@%C%x%�&'        >%@%C%F%        m%x%�&'        {%~%�%�%        {%~%�%�%        �%U&�&�&        �%�%�&�&        �%�%�&�&        �%�%�%�%�%�%        �%�%�%�%        �%�%�%'&�&�&        �%�%�%�%         &'&�&�&        *&-&5&L&        *&-&5&>&        '!'#'&'        O'�'�'�'�' ((((�(�(�(        �'�'�'�'(0(        �'�'�'�'        �'�'`(�(        �'�'�'�'        �'�'�'�'`(�(        `(f(h(k(        �'�'0(`(        �'�'0(`(        0(6(8(;(        �(�(�(�(        �(�(�(�(        �(�(�(�(        �() )')0)})        �)4*+:+        *)*+:+        ****        K*�*�*+:+C+        o*�*�*+:+C+        o*u*x*{*        Z+f+p+}+�+�+        Z+_+b+d+        p+}+�+�+        �+�+�+�+        �+�+�+�+        :,=,C,�,        �,�,�,�,�,�,        �-�/�/0        �-�-�-�-        �-�.�/0        �-.. .        f.i.l.�.        �.�.�.�.        //�/�/        ////        /�/�/�/00        0/6/>/�/�/�/00        S/�/�/�/00        S/Y/\/_/        10i0n0�0        10F0I0L0        �0�0�0�0�01161        �0�0�0�0161        p$r$�$�$�$�$�$�$�$9'@'�(�(})�)�)�)�)�)�)�)C+P+�+�+�+�+�-�-0 0�0�0�0�061@1]1        d2f2i2m2u2�2�2�2        �2�2�2�2        �2�2�2�2�2�2        �2�2�2�2        �2�2�2�2        3333 3:3        D3F3I3M3U3�3�34        `3�3�3�3�3�3�34        �3�3�3�3�3�3        �3�3�3�3        j3�3�3�3�3�3�34        w3�3�34        4G4`4�4        �5�5 6666        (6?6P6g6j6o6�6�6�6�6        (686P6g6�6�6�6�6        ]6g6�6�6        86?6�6�6�6�6        �6�6 7$7(7C7        �6�67 707C7        `7r7�7�7        �7�7�7�7�7�7�7�7        �7�7�7�7        �7	88/8        98J8P8o8p8r8        b8e8k8o8        `1b1p1u1�1�1�1�1�1�1�1�1�1�1�1�1 222&202T2`2�2 3?3@344�4�4�4�4�4�4D5P5�5�5�5�56 6�6�6C7P7�7�7�7�7�7�7/808r8�8�8�8�8�8�8�8�8�8�8 999*90989@9H9P9X9`9l9p9�9�9�9�9�9 :::U:`:e:p:�:        �<�<�<�<        �<�<�<�<        �<�<�<�<        �<�<�<==L=        �<�<�<==L=        �<==L=        �<�<G=L=        �<==G=        e=i=�=�=        i=x=�=�=�=�=        �=�==>B>        �=>>6>;>=>        >6>;>=>        v?y?�?�?�?@        �?�?�?@        �@B B?C        LARAUA�A        �A�A�A�A�BC:C?C        �B�B�BC:C?C        �B�B:C?C        �B�B�BC        �A�A�A�A�B�BC:C        �A�A�B�BC:C        �B�BC:C        �B�BC:C        �A�A�A�A        ���������:�:�:�:�:�:�:�: ;;;B;P;d;p;�;�;�;�;�;�;�;�;�;�;�;�;�; <<<< <(<0<Q<`<�<�<L=P=�=�=B>P>�>�>p?p?@ @h@p@�@�@?C        �C DDDDD        RDTDWD[D_DaDgDmD        �D�D�D�D�D�D�D�D        @CZC`CpCpC�C�C�C�C�C�C�C�C�C�C*D0DKDPD�D�D�D        �D�D�D
FF:G@G�G�G�G�G�G HH        �H�H�H�H�H�H�H I        �H�H�H I        II	II        >I�I�I5J@J~J        HI�I�I0J@J~J        NITIXI[I�I�I�I�I        �I�I�I�I�I�I�I�I        �I�I�I�I        FJOJ`J~J        JJMJ`J~J        OJQJUJWJ        �JK0K<KCK�K        �J�J�K�K        �JKPK�K        �JKPK�K        PKwK�K�K        YKbK�K�K        �K�M�M�M�MP        �K�M�M�M�MP        �K�K�N�N        �N�N�N�N�N�N�N�N        �KLPP        LzL~L M N�N@O�O�OP        @O�O�O P        uLxL~L�L�L�L�L M N�N PP        uLxL�L�L�L�L�L M PP         N*N0N2N5N8N;NBN        CMeMiM�M OOOOO(O        PMeMOO        iM�MO(O        �M�M�N�N        �MNNN        'P+P3P\QpQ�Q�QoRyR�R        ]P�P�R�R�R�R        oPrPvPyP|P�P        �P�P�R�R        �P\QRoRyR�R�R�R        /QOQSQ\Q        3Q7QSQ\Q        RRRRRR        0RgRyR�R        >RBRERNRyR}R�R�R        �Q�Q�Q�Q        �Q�Q�Q�Q        �R�R�R�R�R�R        CSFSSSYS\S_S        |S�S�S�S        OU�U�U^VfVxV        RUZUsVxV        jU�U�UYVfVsV        �U�U�U�U�U�U�U�U        �V�V�V�V        �V�W�WX X@X        WW;X@X        <W�W�W X        <WPWhW�W�W X        <WGWkWW�W�W        GWPW�W X        WXrX�X�X�X�X        �X�X�X�X        �X�X�X�X�X�X        �X�X�X�X        �XvY�Y�Y Z�Z        �X;Y Z0Z        �XY Z0Z        	ZZZZ"Z0Z        �Y�Y�Z�Z        �Y�Y�Z�Z        �Y�Y�Z�Z        �Y�Y�Y�Y        9ZBZiZrZ        �Z�[�[a\p\�\        [![&[3[        ![$[@[D[F[K[M[P[        T[�[�[a\p\�\        �[�[z\�\        �[�[�[�[�[\        �\R]`]�]        �\ ]]]        ] ]`]�]        i]l]s]y]�]�]        �]�]�]u^�^9_        �]�]4_9_        �^�^�^�^�^�^        I_�_�_�_�_�_        m`p`x`�`        �`,a/a1aCaEaOa�a        �`aOa�a        �`�`�`a        Oaha�a�a        �a�a�a�a�a�a        �abb$b        _cbcecyc        �d eeeUele        �f%g(g*g0gpgsgug        �f�fg#g        ggg#g        �g�g�g�g        �g�g�g�g        �g�g�g�g        �g�g�g�g        �g�g�g�g        �g�g�g�g        �gh	hh        0hChGhLh        5hChGhLh        5h8h<h?h        Xhbhehkh        �h�h�h�h        �h�h�h�h        �h�h�h�h        �h�h�h�h        �hiii        �hiii        �h�h�h�h        iiii        Picigili        Uicigili        UiXi\i_i        �i�i�i�i        �i�i�i�i        �i�i�i�i        �i j#j4j�j�j        bj�j�j�j        �j�j�j�j        k`kcktkl$l        �k�k�k�k�k�k        �k�k�k�k        �k�k�k�k        m.m@mZm        BmEmJmWm        cnfnin�n�n�n        cnfninwn        �n�n�n�n        o"o%o9o        ^oaodo�o�o�o        ^oaodogo        �o�o�o�o        �oppp        >pApDpop�p�p        >pApDpGp        �p�p�p�p        �p�p�pq        )q,q/qXq`qzq        )q,q/q2q        bqeqjqwq        �q�q�q�q        	rrr:rPrjr        	rrrr        RrUrZrgr        -s0s3s\sps�s        -s0s3s6s        rsuszs�s        MtPtSt~t�t�t        MtPtStVt        �t�t�t�t        tuwuzu�u�u�u        tuwuzu}u        �u�u�u�u        �v�v�v�v�v�v        �v�v�v�v        �v�v�v�v        BwEwHwXw        �w�w�w�w        �w�w�w�w        �xyy%y        yyy%y        yy%y/y3y8y        hy�y�y�y        �y�y�y�y        �y�y�y�y�y�y        �y�y�yz        o{�{�{�{        �{�{�{�{        �{�{�{�{�{�{         H~H�H I I.I0I~J�J�K�KP P�R S+S0SaSpS�T�T�T�T�T�T@U@UxV�V�V�V@X@X�X�X�Z�Z�\�\�]�]9_@_�_�_�_�_�_�_�_�_�_ `
``` `(`0`:`@`J`P`�`�`�a�a�a�ab�bMcPc�c�c�d�d�e�e�f�fyg�g�g�g�g�gLhPh�h�hiilipi�i�ikkGlPl�m�moo�o�o�p�p�q�q�r�r�s�s�t�t v v w w]w`w�w�w�w�wx x{x�x�x�x8y@yOyPy�y�y�y�yEzPz�z�z�z�z1{@{O{P{�{�{�{�{�{�{8|@|G|P|b|        �|�|�|�|        �|�|�|�|        �|�|�|�|        0}4}8}F}        0}4}8}:}        P}T}X}Z}        4~8~<~f~        t~x~|~�~        ����        ����        ����        ����        ����        ����        ����        ����        ����        0�4�8�<�        ��������        ��������        ��� �	�P�a�        ��� ��        ��� ��        �,�C�I�        '�+�/�F�P��        '�+�/�1�3�6�        '�+�/�1�        C�L�T�]�p���        C�G�T�Y�        C�G�T�V�        p�s�u�x�z�������        ��������Ѓ������        ������������        ��������        Ѓ����        q�u�z�������        q�u�z�|�����        q�u�z�|�        ��	�#�%�        �����������������        ������������        ��������        g�k�w�|�~���        g�k�w�y�        #�'�/�4�        #�'�/�1�        w�{�������χ҇ԇ��        w�{���������        w�{�����        A�E�J�X�`���        A�E�J�L�Q�T�        A�E�J�L�        ������������        ��������        ������������        ��������        ��������        ӈ׈߈��+�        ӈ׈߈��+�        ӈ׈߈�        ӈ׈߈�        �����        ������        �����        ����        7�;�G�������        7�;�G�P�����        7�;�G�L�        7�;�G�I�        P�]�����        o�}�����        ǉˉω��        ǉˉωԉ        ǉˉωщ        ������        ���Q�Y�j�        ����Y�j�        ����        ����        ?�A�L�Q�        u�y�������ʊ        u�y�������ʊ        u�y�����        u�y�����        ��������        ��������        |�ԋً�        �����        �?�P�p�        ��"�7�P�`�        7�?�`�p�        Ԍڌ܌ߌ         �-�.�3�         �&�(�+�        M�U�`���        `�f�h�k�        ������$�0�����C�        ��������        ��������        �����0�`��C�        ύӍٍۍ        Ӎ֍ۍ����� �        ֍ٍ��        �� �C�         �&�(�+�        ����        F�`� � �        |������        �$�����        ѐ���        ����ő֑        ���
���        ����        (�,�0�6�D�q�        �������        ��ؒ���        ��ؒ���        D�I�M�]�        ��������        ˓�����        ˓ϓғԓ        *�.�N�_�        ��������        ����	�        ����	�        �!�'�*�        !�'�*�0���ƕ        �����        �����        �����        ��+�<�        ǖԖ��        Ԗ��!�        �� ��        �A�P����������        ,�A���������        ��������        T���З�        X�f���        n���З�        ������З        W�[�k�y�        W�[�k�p�        W�[�k�m�        y�}�����        ��"�3�        ��"�3�        K�N�T�W�        g���ę�        ������������ʙ͙        ����͙љ        ����ęʙљ�        �4�P�t�        "�$�'�*�        $�'�*�2�P�t�        P�V�X�[�        ߚ'�@�p�        �'�@�p�        ��S�`�         �'�`�p�        ��������0�A�        ��������        ��������        ���� �0�        ؛�� �        ��� �0�        g������        g�{���        g�i�n�q�        ����ǜМ���        ����М��        ���� ��        ����M�        ��ǝ@�M�        ��������        ��� �0�        ���0�@�        `�r�����������Ǟ        `�b�g�j�        b�g�j�l���Ǟ        ��/�@�N�        (�/�@�N�        k�������        ��������        ߟ���        #�)�,�/�        )�,�/�;�P�c�p�x�        3�;�p�x�        ;�A�c�i�        ��������        �������        ����������        ���� ��        �������        ��ƠȠˠ        2�j�x���        �����        �2�?�\�        o���âТӢآ��        v�x�~���        ��������âТ        ������        �� �s�x�         �V�c�p�����        #�%�+�-�        3�9�>�N�c�p�        N�V�����        ��������        ����ӣ�        ������ǣ         �	��/�        5�9�A�C�        S�W�r���        ������        ������ �0�        äŤˤͤ        Ӥ٤ޤ���        ��� �0�        7�=�C�J�        i�l�r���Х���������        i�l�r��̦ߦ        i�l�r�w�        i�l�r�t�        ������̦        �P�ߦ��        ���P�        ����        %�+�-�0�        P����������        c�f�l�n�        i�l�r������        7�;�K�]�        7�;�K�P�        7�;�K�M�        ]�a�����        ԧاܧާ        ������        ������        ������        l�p�t�v�        ��������        ĨȨ̨ݨ        ĨȨ̨Ψ        ������        � �$�&�        ��������        p|w|�|�|�|�|�|�|�|�|�|�| }+}0}G}P}m}p}�}�}�}�}#~0~f~p~�~�~�~�~&09@FP[`s�������������"�0�?�@�J�P�Z�`�f�p�z�����������ǀЀ׀�����a�p�����ɁЁ����� ���� ������5�@������ �>�@�e�p�����*�0�N�P�u��������� �� �E�P�^�`�͆І���� �e�p������5�@�����ÈЈ+�0������� �j�p�ʊЊۊ������� ���� �,�0�S�`�h�p����p�p�������������ŌЌ��3�@�����C�P������������� � �S�`�����������0�0�c�p�����֑��� �x�����2�@�d�p������� �_�`�����������ƕЕ��<�@�a�p�u�������!�0�C�P�����՘���� �3�@�X�`���t���Кp�p�u���A�P�� �%�0�Q�`�e�p�����M�P�ǞО��R�`�ğП� �x������ �������\�`���������/�0�����0�0�T�`��� �"�0�����ȧЧ��� �S�`���������ݨ���5�@�w�����������ЩЩ����0�        4�:�<�?�        M�P�S�]�p�|�        M�P�S�V�        V�]�p�|�        ݫ��� ��        ݫ���        �� ��        m�p�s�}�����        m�p�s�v�        v�}�����        �� ��� �,�        �� ���        �� �,�        ������������        ��������        ��������        O�R�U�_�r�~�        O�R�U�X�        X�_�r�~�        ݮ��� ��        ݮ���        �� ��        m�p�s�}�����        m�p�s�v�        v�}�����        �� ��� �,�        �� ���        �� �,�        ������������        ��������        ��������        �-�@�J�        � �#�&�         �#�&�-�@�J�        |�����������űѱ���        ��������űѱ        ��������        ����űѱ        �	��G�J�S�^�d�i�u�����        7�:�=�G�i�u�        7�:�=�@�        @�G�i�u�        0�T�`������������ �����6�@�ƬЬV�`�������6�@�ƯЯV�`���]�`��� �����òв�        ����������ϳ        ��������        ������ϳ        ��������        ����         �/�0�Q�`��        �#�0�f�p�ŵ͵c�        M�P�V� �0�f�p���͵c�        M�P�V���0�E�p���͵�        e�t���        t�����˴p���͵�        t���v�x�{���͵�        v�x�{���͵ٵ        v�x�{���        ��������        ����´˴        ����N�U�        K�N�S�f�        ���;�        �c�        p�v���������        ������з        ���зܷ        ��зܷ        2�z�зܷ        H�Q�W�Y�        ��'�7�d�������        '�7�d��������&�.�_�        '�I�d�p�����        r�7������&�.�����_�        r�}���ظ�7������&�.�����_�        ����P���7�.�����_�        ��������7����H�_�        ��»�"�        ��e�j��1�        ����        �"�&�*�.�2�        �"�&�*�        �"�&�(�        6�E���        ��� �������        ��� �p�����        ��O�X�� �p�����        {�}����        }������        ��϶ж� ���_�`���        ����        ��������        �4�@�]�p�~�        ���"�        ������������        ���� �~����� ��         �"�0�2�@�F�P�V�`�e�p�u�����������������        !�>�P�U�        ���������������� ���Y�        ��������        7�;�=�S�        ����
�        -�G�x�������        -�G�x�������        `�������������� �����
����        �����������        �O�P�^�`�l�p�~�����������������        ����������	�        ��	��� �,�        5�V�Y�\�`���        ��� �]�        0���������]�`���        �����������        �������        ���         �&�0�?�@�a�        p������        ��������        ��������������        	��1�3�        �/�3�;�        ��������        ����        ����3�@�c�p���        ?�[�b�v�        �������        ����������� ������        <�����A�a���        <�A�H�M�        A�H�M�����������        ��A�a�o�        ���        ��������        ����        �����������        Q�[�n�p�w����������        <�C��������        6�O�R�W�����        O�R�W�j�        j�~���5�        ~���5�[���        n�����9�        ����9�_�����        ��� ���        ������        ������ �        ������ �        #�,�P�\�        i�o�r�����q�        i�o�r�z�0�:�        z�����0�:�q�        z�������        ������ ��0�        ������ ���        ������ �        �����0�        ����        S�Y�[�^�         �H�P�%�0�W�`���������� �\�`�q�        ������������        ��������        ��������        ��������        ������������ �P�        a�g�o�t�y�|�        ������        P�S�`� � �����������"�0�q�        ��������        ��������        ��������        d�y�����        0�L�N�Q�        �����        ������������ �%�0�7�@�O�P�]�`����������� �����A�        P�D�P�������        ���%�        �������        ������        �������        
�T�[��� ���        v��� �[�p���        v����������        v������        ����������������        �������� ���@�        ���� ���@�        ���� �����@�         ���� �@�        ����@�[�p�y�        ����@�I�        ����p�y�        J�T�[�`�        ������_�p�����;�        ��_�p�����;�        ������[�p�����������        ������        �:�=�@�        G�J�R�U�X�[�        G�J�R�U�        w�z���������        w�z�����        ��������        �������-�        ��������        ���������        F�I�O���������n�        a���������n�        a�c�j�������        u�|�����        |�������        ��������        ���F�K�P�`�        �	���        &�)�.�8�K�P�        u�x�������s�        �������        �#�K�P�U�e�        ���#�        .�1�6�@�P�U�        ��������        ����������&�0���        ����0�<�        ������������        d�������        o�r�u���        ���&�        �������� ���        ��0�<�        ��$�&�        T�t���������        _�b�e�t�        �����������        ��������        �����������        �������         �,�[�l�����         �,�e�l�        [�e�����        �0�]�b�g�w�        ��!�0�        ;�>�C�M�b�g�        ��������        �������        �������        ��������        ��"�� ��        ?��� ���        S�_���������        v���p���        ���� �p�        ���� �,�        ����@�p�        ������������        �������        ��������        �����        +�@�`���        2�6�����        6�@�`���        ������������ ���        ���� ���        ���� ��        ���� ��        ���2�        2�R�}�������        =�@�C�R�        ]�`�e�o�����        �����������$���        �������$�P�\���        ��������        �	���        /�2�5�?�����        \�������        g�j�m���        �������������)���        �����)���        ������        )�I�t�y�~���        4�7�:�I�        T�W�\�f�y�~�        ������ ��� ���        �� ��� ���        �� ��� �@�        ���� �,�        ������ �        B�E�J�d�        d�����������        o�r�u���        ������������        ��s�����        !�s�����        !�`�����        2�P�����        2�>�����        @�B�E�H�        `�c�f�i�        ������������        ��������        ������������        
�Y�`����������        =�Y�`����������        =�Y�`���        N�Y�`�n�        ��������        ��������        �����������        ��������        ������������        $�'�-�_�p�u��������        ?�_������������        ��������        �����������        ��������        ������������        %�(�1�]�s������        s�������        �������� ��        ��������        ���������� �        ,�e�v�9�        X�e�v�9�        v�������        ��������        �������+�        ��������        ���������        R�����Y�        ~�����Y�        ��������        ��������        ���1�6�;�K�        �������        ���#�6�;�        v�y�|���	�_ b e p �         v�y�����        ��������� �         ��������        ����"�%�(�/�1�0         ����,�/�1�0         ����,�/�1�@�H�0         ,�/�1�@�P�0         	�"�%�(�0 D p |         	��0 <         �"�%�(�p |         �"�%�(�        J M R _ b e         � � � �  0�         0�         0A        0<        CFKb        b�����        mps�        ������        .<Pip�        .4P]bfp�        P]p�        SW��        W]p�        ����        ����        48:A        TXZa        vy���        ����        ����        ��        ���        ;fkp�        &),;        FINXkp        ��� 7A�        � 7A�        ���AK        ��AK        "%*7        Kk����        VY\k        vy~���        ���>Pgq�        �>Pgq�        ���7q{        q{        RUZg        {�����        ����        ������        	n���        !n���        !#*g��        7;��        ����        ����         ����        �����         69?����N	        Q����N	        QSZ���        gk��        ����        ��&	+	0	@	        ����        					+	0	        f	i	o	�	�	�	
~
        �	�	�	�	
~
        �	�	�	�	

        �	�	

        �	�	�	�	        
+
V
[
`
p
        


+
        6
9
>
H
[
`
        �
�
�
�
'1�        �
�
'1�        �
�
�
�
1;        �
�
1;        '        ;[����        FIL[        finx��        ���.@Wa�        �.@Wa�        ���'ak        ��ak        BEJW        k�����        vy|�        ������        ���^p��        ^p��        W��        '+��        ruz�        �����         ����        ������        &)/����>        A����>        ACJ���        W[��        ����        �� 0        ����        ���         VY_����n        q����n        qsz���        ����        ����        �FKP`        	        &).8KP        ������������ �2�@�O�P����� � �6�@�F�P�k�p���������� �R�`���������;�@�n�p�s������������������ ����������������������� �� �� �� �9�@�Y�`�h�p�� � �����  ������'0BPbp�����������  %0N	P	U	`	~
�
�
�
�������� >@EPnpu        ���	        !0Y^`        !0U        ����        ���0\^a        ���        E\^a        ����������        ����        9�������        ?�����        ����        BDKknp��        cp���}����� '0����4@��� `        `{        ������        ����        ����        ����        "-@`        "%        %-@`        @FHK        �������� !0?@ap�������``op�������� ;@z�������� :@]`}��        �S`�        �s��        ����        �����DP[`cps        � h!        p!v!�!�!�!�!        �!�!�!�!�!>"        A"C"G"�"�"�"        �"�"�"Y#p#�#        #;#>#C#        �!>"@"�"�"�#        b$�$�$�$ %%%%0%�%        s$�$�$�$0%�%        �$�$0%P%        �%�%�%�%        �$�$%%        �$ %% %        �$�$%%        �$ %% %        �$�$�$�$        �%�%&#&0&H&`&s&�&�&�&�&        �%�% &#&E&H&`&s&�&�&        �&�&�&�&        �&�&�&+'        �#�#�#�#�#$$$ $A$P$�%�%�&�&4'        �(�(�(�(�(�(        @'F'P'V'`'t'�'�'�'�'�'�'�'�'�'�'�'( (I(P(_(`(�(�(�(�(�( )))) )&)0)z)���        �)�)�)�)        �)�)�)�)�)�)        $   '   )   >             :  F  �  �  �             ?  P  [          �  �  t            �  �  t            �  �  �            �  �  �  �  �  �          �  �  �  �  �  �          �  f  p  t          �    !  P          �  �  �  �  �  �  �  �          W  }  �  �          �    0  �  �  �          2  r  �  �          	  0	  @	  c	  p	  �	           
  1
  3
  9
  ;
  A
  D
  �
          �
  �
  �
  �
  �
  �
  �
  �
  �
  @          �  P  �+  ,  �,   -  �-  �-  2  C2  �2  �2          �  �  �  �  �+  ,               #  *  �+  �+          X  �  /  2  4  p  u&  �&  3(  �(  )   )   -  #-  �1  �1          X  �  3(  �(  )   )  �1  �1          X  [  3(  e(          e(  �(  �1  �1          h  d  �!  �!  $  0$  �1  �1                   #  )  ,  d          �  �  �  �  �  �  �  P          P  a  g  m  s  x  {  �          �  �  �  �  �  �  �  P          P  a  g  m  s  x  {  �          �  �     �             %  (  1  3  9  B  G  K  �          �  �  �  �  �  �  �            	  1  v+  �+          T  �  g'  3(   )  )  o,  �,  �0  �0  /1  �1  �1  2          �'  �'  �'  �'  �'  �'  �'  �'  }1  �1          �'  3(  R1  }1           )  =)  @)  G)  I)  P)  �0  �0          U)  )  �0  �0          �  �  �  �  �  �  �  #          #  �  �!  _"  �&   '  F0  q0          @  Q  W  ]  c  h  k  �           "  "  "  "  "  $"  '"  _"          �  �  �  �  �  �  �  #          E  �  �#  $  )  �)          p  �  �  �  �  �  �  �          �  �  �  �  �  �  �  �            )  �-  �-            �  �0  /1          �  7  �*  +  0  40          �  v  0$  �%  F.  {.            !  '  -  3  8  ;  v          0$  A$  G$  M$  O$  T$  W$  �$          �$  �$  �$  %  %  	%  %  %  %  O%          O%  �%  F.  {.          v  �  �)  *          �  Y  t-  �-  p/  �/          �  �  �  �  �  �  �  �          �              S          {  �  +  D+          �  �  �  �  �  �  �              �  {.  p/  �/  0  �1  �1          �.  /  �1  �1          �  �  �  �  �  �  �  /          p  �  $  $  #-  `-          ]   �   �)  �)  �1  �1          �   �   �   �   �   �   �   !          �"  �"  D+  v+          0#  A#  G#  M#  O#  T#  W#  �#          �%  �%  �%  �%  �%  �%  �%  �%          &  !&  #&  )&  /&  4&  7&  u&           '  '  '  '  '  $'  ''  g'          *  �*  `-  t-  �1  �1  C2  �2          0*  S*  �*  �*          {*  �*  `-  t-  �1  �1  C2  �2          �*  �*  �*  �*  �*  �*  `-  t-          X2  b2  d2  �2           3  3   3  '3  �8  9          P3  a3  g3  m3  s3  x3  {3  �3          �3  �3  �3  �3  4  4  4  `4          `4  q4  w4  }4  �4  �4  �4  �4          �4  �4  �4  �4  5  5  5  P5          P5  v5  9  F9          v5  �5  �8  �8          �5  �5  x9  �9          �5  �5  �5  �5  �5  6  6  P6          Y6  �6  �9  :          �6  �6  �6  �6  �6  �6  �6  @7          @7  Q7  W7  ]7  c7  h7  k7  �7          �7  �7  �9  �9           8  8  8  8  #8  (8  +8  p8          |8  �8  F9  x9          �:  �;  �;  �=          0;  A;  G;  M;  O;  T;  X;  �;          �;  �;  �;  +<          +<  <<  B<  H<  J<  O<  S<  �<          �<  �<  �<  1=          �<  �<  �<  �<  �<  �<  �<  �<  �<  1=          1=  B=  H=  N=  P=  V=  Z=  �=          �=  �=  p>  p?  @  0@          �>  �>  �>  �>  �>  �>  �>   ?          �=  >  0@  b@          >  +>  �?  �?  �?  �?          �?  �?  �?  �?          @>  _>  p?  �?          �@  A  A  'A  dC  �C          A  A  'A  dA  /B  GB  PB  WB          �A  �A  �B  �B  �B  �B  �B  �B          �B  �B  �B  �B          �A  �A  �A  �A   C  2C          rB  �B  �B  �B  2C  dC           D  �D  �D  �E          3D  GD  ID  PD  �D  �D          oD  �D  �D   E           E  PE  wE  �E          PE  wE  �E  �E          F  !F  #F  )F  +F  0F  3F  pF          �F  �F  �F  �F  8G  �G          �F  �F  �G  �G          �G  tH  �H   I          �H  �H  �H  �H          pI  �J   K   L  $L  *L  @L  �M  �M  �f          pI  �I  �I  �J   K   L  @L  �M  �M  �f          �I  �I  �I  �I  �I  �J  �J  �J  K   L  @L  �M  �M  �f          �I  �J  �J  �J  K   L  @L  �M  �M  �f          -J  �J  K  �K  �L  �L   M  �M  �M  �M  4N  8O  YO  rO  �O  xe  �e  �f          aJ  �J  �M  �M  4N  �N          XK  �K  �N  8O  �O  �Q  �R  �R  �R  V  �V  �Z  �Z  @]  P^  _  _  p_  ~_  �_  �`  �a  �a  �c  �c  �c  �c  Od  �d  xe  �e  �e  �e  �e  0f  af  f  �f          �O  :P  SS  �S  T  jT  �U  �U  �U  �U  X  kX  �Z  \  $\  �\  �^  _  �`  a  Da  �a  b  Pb  sb  �b  �b  �b  Mc  �c  �d  e  �e  �e  f  �f  �f  �f          �O  &P  �U  �U  �Z  \  $\  �\  Da  �a  b  Pb  sb  �b  �b  �b  ^c  �c  �d  e  �e  �e  f  �f  �f  �f          P  &P  Da  �a  �e  �e  �f  �f          �U  �U  �Z  �[  sb  �b  �b  �b          $\  �\  b  Pb  ^c  �c  �d  e          $\  7\  b  *b          &P  :P  �`  a  �f  �f          T  jT  �^  _          .T  IT  KT  OT          )X  UX  Mc  ^c          :P  �P  �S  �S  �T  U  ]U  �U  �U  V  �V  X  �Z  �Z  \  $\  �\  �\  P^  �^  _  p_  ~_  �_  �a  �a  �a  b  �b  �b  �c  �c  .d  Od  e  xe  �e  �e  >f  af          �P  �P  �U  V  �V  �W  P^  �^  _  p_  �a  �a  �a  b  �c  �c  e  xe  �e  �e  >f  af          �P  �P  _  p_  �a  �a  �e  �e          �U  V  �V  tW  �a  b  e  )e          P^  �^  )e  xe  >f  af          P^  c^  Je  `e          �P  �P  �\  �\  .d  Od          �T  U  ~_  �_  �b  �b          �T  �T  �T  �T          �W  X  �e  �e          �P  �Q  �R  SS  jT  �T  U  ]U  �U  �U  X  X  kX  �Z  �Z  �Z  �\  @]  a  Da  �a  �a  Pb  sb  �b  Mc  �c  .d  �e  �e  0f  >f  �f  �f          BQ  �Q  �U  �U  kX  vY  �Y  �Z  �\  @]  Pb  sb  �b  Mc  �c  .d  �e  �e          rQ  �Q  �\  @]  6c  Mc  �e  �e          �X  OY  �b  6c          �Y  �Z  Pb  sb  �c  .d          �Y  Z  �c  d          U  ]U  �U  �U  �a  �a          vY  �Y  0f  >f          a  Da  �f  �f          M  �M  �Q  �R  �R  �R  V  �V  �Z  �Z  @]  P^  _  _  p_  ~_  �_  �`  �a  �a  �c  �c  �c  �c  Od  �d  �e  �e  �e  0f  af  f          M  +M  �Q  �Q          �Q  �R  �R  �R  V  �V  �Z  �Z  @]  P^  _  _  p_  ~_  �_  �`  �a  �a  �c  �c  �c  �c  Od  �d  �e  �e  �e  0f  af  f          8R  �R  �Z  �Z  @]  P^  �_  �`  �a  �a  �c  �c  �c  �c  Od  �d  �e  �e          hR  �R  vd  �d  �d  �d  �e  �e          �]  P^  �a  �a  �d  �d          �_  �`  �c  �c  �c  �c          �_  `  �c  �c          V  TV  �Z  �Z          �_  �_  �e  �e          �J  �J  �L   M          �K   L  N  4N          �L  �L  rO  �O          �L  �L  �M  N  8O  YO           g  Gh  Kh  Qh  `h  %i  0i  �m  �m  n           g  h  `h  #i  0i  @i  Bi  Ei  Pi  �m  �m  n          *g  	h  `h   i  0i  @i  Pi  �m  �m  n          vg  �g  �h   i  `i  �j   k   l  `l   m   m  nm  �m  �m          �g  �g  `l  �l  �m  �m  �m  �m          �i  �j  �l  �l  �m  �m          2k   l   m  nm          2k  Ek  @m  Vm          �g  	h  �j  �j          �h  �h  �j   k          �j  �j   m   m           l  `l  nm  �m          Sn  ]n  `n  �n   o  �p  �p  �s  �s  #�          `n  �n   o  }p  �p  �s  �s  #�          �n  �n  �t  �t          6o  Pp  �p  �q  �q  �q  r  �s  �s  t  Gt  ct  �t  �t  �t  �w  �w  ؍  �  #�          eo  Pp  Gt  ct  �t  �t  �t  Gu  �w  Rx  zz  �z  �z  �z  �z  |  }  �}  �~  �~  �  4�  ��  ߀  ��  �  ��  щ  j�  ��  ؊  ��  �  l�  �  �  �  $�  a�  ��          uo  p  �t  Gu  �w  Rx  zz  �z  �z  �z  �z  |  }  �}  �~  �~  �  4�  ��  ߀  ��  �  ��  щ  j�  ��  ؊  ��  �  l�  �  �  �  $�  a�  ��          �o  p  �z  �z  �z  |  }  �}  �  4�  ��  �  ��  щ  x�  ��  �  l�  �  �  �  $�  a�  ��          �o  p  ��  �  �  �  �  $�          B{  |  <�  ^�  a�  ��          9}  �}  ��  щ  �  <�  ^�  l�  �  �          9}  H}  �  $�          
x  Rx  zz  �z          �~  �~  j�  x�          ��  ߀  ؊  ��          q  �q  Zu  pw   y  y  �y  zz  �z  �z  |  }  �}  �~  �~  �~  4�  b�  ��  ��  �  _�  ��  ��  ��  s�  ��  ��  щ  �  ��  Ȋ  ��  �  l�  �  �  ��  ��  ��  �  �  $�  a�  ��  Ԏ  ��  �  /�  B�  P�  ��  ��  #�          Zu  v  *z  zz  |  L|  �|  }  �~  �~  �  �  ~�  ��  ��  ��  �  $�  щ  �  ͋  �  l�  w�  �  ��  P�  ��  T�  ��  Đ  ʐ  ѐ  ��          �u  v  �~  �~  ��  ��  ͋  �  l�  w�  <�  ��  ^�  ��  T�  ��  Đ  ʐ  ѐ  ��          �u  v  ͋  �  l�  w�  T�  k�          �  ��  k�  ��  Đ  ʐ  ѐ  ��          �  ��  <�  ��  ^�  ��          �  ��  O�  e�          �|  }  �~  �~          �  $�  P�  ^�          щ  �  �  <�          v  �v  �y  �y  �|  �|  E~  �~  K�  b�  ��  ��  ��  �  `�  s�  ��  ��  ��  Ȋ  ��  D�  ��  ��  �  �  $�  /�  ��  �  ��  �  %�  )�  .�  T�  ��  Đ  ʐ  ѐ  ��  ��          ^v  �v  [�  b�  `�  s�  ��  ��  ��  D�  ��  ��  $�  /�  ��  �  ��  �  %�  )�  .�  T�  ��  Đ          �v  �v  ��  D�  $�  /�  ��  �          ��  N�  ۏ  ��  %�  )�  .�  T�          �  ��  ��  ۏ  ��  �  ��  Đ          �  �  ��  Ï          O~  �~  K�  [�  ʐ  ѐ          ��  �  �  �          ��  Ȋ  �  �          �v  pw  �y  *z  L|  �|  �}  E~  4�  K�  ��  ��  �  _�  ��  ~�  ��  ��  $�  `�  D�  ͋  w�  �  /�  a�  ��  Ԏ  /�  B�  ��  ��  �  %�  )�  .�  ��  #�          w  pw  D�  K�  �  _�  ��  ~�  D�  ��  w�  �  /�  a�  ��  Ԏ  /�  B�          <w  pw  D�  ��  w�  ��  ��  Ԏ          l�  8�  /�  Q�  ��  ��          ��  ~�  ��  �  /�  B�          ��  у  ��  ��          �}  E~  4�  D�  �  %�          $�  `�  ��  ��          ��  ͋  ��  #�          Rr  �s  Gu  Zu  pw  �w  Rx   y  y  �y  �z  �z  �~  �  b�  ��  ߀  ��  _�  ��  ��  ��  s�  ��  �  j�  Ȋ  ؊  ��  ��  ��  ؍  Ԏ  ��  �  /�  B�  P�  ��  ��          Rr  dr  pw  �w          dr  s  Rx  �x  �x   y  y  ay  �z  �z  �~  �  b�  ��  ߀  ��  _�  ��  ��  ��  s�  ��  �  j�  Ȋ  ؊  ��  ��  ��  ؍  Ԏ  ��  �  /�  B�  P�  ��  ��          �r  s  �z  �z    �  ߀  ��  ��  ��  s�  ��  �  j�  Ȋ  ؊  ��  ��  ��  ؍  �  /�  B�  P�  ��  ��          �r  s  s�  ��  ��  ��  ��  ��          Q  �  $�  D�  ��  ؍          ��  ��  �  $�  D�  j�  �  /�  B�  P�          ��  �  D�  Z�          y  ay  �z  �z          /y  Gy  Iy  My          _�  ��  Ԏ  ��          Zp  }p  �s  �s          �p  �p  �q  �q          t  Gt  �w  �w          t�  #�  &�  )�  C�  ��  Л  �  6�  ��  ��  Ǟ  �  �  v�  �  |�  ��  ʢ  ڢ  �  ��  ��  �  �  ��  �   �  C�  d�          ~�  #�  C�  ��  Л  �  6�  ��  ��  Ǟ  �  �  v�  �  |�  ��  ʢ  ڢ  �  ��  ��  �  �  ��  �   �  C�  d�          ˑ  #�  ��  Ǟ  �  �  Ƞ  �  ʢ  ڢ  �  ��  ��  �  �   �          ��  #�  ��  �  ��  ţ  �   �          3�  �  �  L�  ţ  �          �  ��  �  �  L�  ��          �  ��  L�  b�          @�  ��  ��  ��          v�  ��  �  ��          |�  ��  C�  d�          p�    В   �          p�  Г  �  8�  Y�   �  s�  C�    Л  �  6�  ��  ��  Ǟ  �  �  v�  �  |�  ��  ʢ  ڢ  �  ��  ��  �  �  ��  �   �  C�          Y�  �  
�  �  s�  C�    Л  �  !�  (�  6�  ��  ��  Ǟ  �  �  v�  �  |�  ��  ʢ  ڢ  �  ��  ��  �  �  ��  �   �  C�          c�  �  s�  ��  ��  C�    Л  �  �  (�  6�  ��  ��  Ǟ  �  �  v�  �  |�  ��  ʢ  ڢ  �  ��  ��  �  �  ��  �   �  C�          ��  �  ��  m�  ��  ��  0�  v�  �  "�  C�  |�  ڢ  �  ��  ��  �  �  ��  �   �  C�          ޙ  �  0�  v�  �  �  ��  �          ��  m�  �  �  ��  ��          �  ��  C�  |�  ڢ  �   �  C�          �  ��  C�  Y�          }�  ��  Ǟ  �          ��  C�  �  �          m�  ��  ��  ʢ          �  0�  "�  C�          P�  ��  8�  Y�          ��  ��   �  g�  ��            �  ��  �  !�  $�  -�          �  ��  �  �          b�  �  ��  ��          w�  z�  ��  	�          y�  ��  ��  ��          y�  ��  ��  ��          ��  ��  ��  ��  ��  ��          �  6�  ��  Χ          4�  6�  ��  Χ          ;�  ��  ��  ��          �  ��  ��  ��  ��  ��          ��  ߨ  �  �          ��  ��  ��  ��          ��   �  3�  5�  ��  ݫ          ܩ   �  ��  0�  ī  ˫          ��  ��  Ū  �  ī  ˫          ��  ��  Ū  ڪ          O�  U�  [�  ��          O�  U�  [�  m�          �  %�  P�  ��  ��  �  &�  5�  <�  k�          b�  ��  ��  �  &�  5�          %�  '�  i�  0�  @�  P�  �  &�  5�  <�  k�  ��          ��  ��  ��   �  @�  P�          ��  ��  �  �          ��  ��  Э  @�          Ѱ  `�  c�  e�  ��  ��  �  �  P�  s�          �  0�  ��  ��  �  �  P�  s�          ��  ��  P�  s�          p�  ��  ��  �   �  P�  s�  Զ          ��  ��  s�  P�  @�  ��  ��  Զ          Y�  w�  }�  ��          �  7�  ��  й  к   �          o�  з  p�  `�  ��  ��  �  к  P�  �  �  ~�  ��  	�          ��  з  u�  �  ��  	�          ��  `�  0�  ~�  ��  ��  ��  ݼ          ��  и  P�  f�          �  к  �  0�  ��  ��  ݼ  ��          ַ  0�  @�  P�          `�  ��  �  �           �  @�  ~�  ��          ��  ��  ��  ��  Ľ  ڽ  �  �  
�  �   �  *�          ��  Ľ  ڽ  �  �  
�  �   �  *�  ſ  �  �  �  �  !�  d�          Y�  ]�  f�  ��  G�  d�          �  ��  ��  o�  ��  ��          ��  ��  o�  ��  ��  ��  ��  ��          ��  ��  ��  ��          �  �  <�  G�          ��  �  �  �   �  G�          ��  ��  ��  ��             
      H   `   �   �   �   �   �     9          q   �   2  9             @   P   |   �   �   �   X  `  u          ~   �   �   �     -          �   �   �     @  +
          B  G  J  L  T  }          �  �  $  �  E	  s	  x	  
          �  �  .  �  E	  j	  x	  
          �  �  .  j  �	  �	  �	  
          j  �  E	  j	  x	  �	  �	  �	          �  �  
  +
          �  �  �  �          .  2  8  Y          �  �    +          �
  �
  �
  �
          �
  �
  �
       �     �  �  �  �  T  p  �  �  &     �  �  �          �  �  0  �  p  �  �  &     p          �  �  3  5  9  y  �  �  p  �  �  �  �  &     p          �  �  t  y  �  �  p  �  �  �  �  &  @  P          �  �              3  5  9  t     @  P  p          �  �  \  �  &  Y  �     �  �          �  �  \  �  &  P  �     �  �          �  �  \  �  �  �          �  �  �  �  &  P  �     �  �          �  �  �  �          �    �  �  �  �          0  G  N  P          a  g  l  p              &  �  �  �          �  0  :  �  �  �  �  '  >  �          �  �  �  �  �  0  :  �  �  �  �  '  >  �          �  �  :  M  �       '          �  �  �  0  M  �  �  �       >  �          @  W  �  �          �                 �  �  o  r  t  {  }  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �  �    	      '  )  7  9  >          �                4  b  �  �          S  W  `  y          �  �  �  �  R  u          R  Z  ^  u          <  X  @  G          L  P  T  p          p  t  z  �          �    0  @          �    0  @          �    0  @          �  �  p  �  �  �          p  t  x  �  �  �          �  '  @  D          �  '  @  D          �  '  @  D          p  �  �  �               �  �  �  �          @  �  �  �          0   f   �   �   !  `!  �!  �!          X   f   !   !          f   p   w   ~   �   �           �   �   �   �           �   �   `!  f!          �$  �$  %  %          #%  )%  B%  O%          i%  �%  �%  �%          '&  D&  J&  M&          �&  '  '  '          �'  �'  �'  �'          P(  �(  �(  �(          �   �   �   �           �  �  �  �          �  �  �  �          �  �  �  �  �  �  �  �          �  �  |  ~  �  �          *  .  6  :  P  n  ~            *  .  6  :  �            n  t              Z  ^  f  j  �  �  �  _	  b	  d	          Z  ^  f  j  �  M	          �	  �	  �	  �	          �	  �	  �	  �	          N
  �
  �  �  8  C          a
  �
  �  �  8  C          �
  4  �  `  @       8  C  ~                          '  a  p  y          a  `  @  �  �  �  C  p  y  ~          �  `  @  �  �  �  [  p          �  �    `  @  L          �  �                   #  �              5  @  G  I          |  @               �  �  �  @                     K          �  �  �             .symtab .strtab .shstrtab .init .text .fini .rodata .eh_frame .gcc_except_table .tbss .ctors .dtors .jcr .got.plt .data .bss .comment .debug_aranges .debug_info .debug_abbrev .debug_line .debug_str .debug_loc .debug_ranges                                                    ���                     !         ���   bh                '         �i 
                  -         @�@i T         @       5         ��	�u �                ?         � �                 Q        D�                   W         D�                    ^         0D0�                   e         8D8�                   j         <D<�                  s         `D`� x                   y          Eش H&          @       ~      0       ش                  �              �  +                 �              �� �,                �              � �v                �              U� �S                �      0       � �               �              �� �#                �              �" ��                              "�# �                                �# �    �1        	              �3' �Q                                    ��          ��          �          @�          ��	                    D          D          0D     	     8D     
     <D          `D           E                                                                                                                                  ��   @�         A�      -   B�      >   C�      U   D�      j   H�      v   L�      �   P�      �   T�      �   X�      �   \�      �   `�      �   d�      �   h�        l�      %  p�      M  t�      ~  x�      �  ��      �  ��      �  ��      �  ��      �  ��        ��      B  ��      Z  ��      q  ��      �  ��      �  ��      �  ��      �  ��      
  ��      5  ��      d  ��      �  ��      �  ��      �  ��      �  ��      �  ��      �  ��        ��        ��      "  ��      0  ��      D  ��      X  ��      o  ��      }  ��      �  ��      �  ��      �   �      �  �      �  �      �  �      �  �        �        �      +  �      @   �      U  $�      i  (�      x  ,�      �  0�      �  4�      �  8�      �  <�      �  @�      �  D�        H�      1  L�      Q  P�      m  T�      �  X�      �  \�      �  `�      �  d�        h�        l�      <  p�      R  t�      j  x�      �  |�      �  ��      �  ��      �  ��      �  ��        ��      9  ��      X  ��      w  ��      �  ��      �  ��      �  ��      �  ��      	  ��      E	  ��      p	  ��      �	  ��      �	  ��      �	  D      �	  0D     	 �	  ��	      �	  8D     
 
  ��      
   �      /
  `�      E
   E     T
  E     b
  ��      n
  E                 ��   �	         �	      -   �	      >   �	      U   �	      j   �	      v   �	      �    �	      �   $�	      �   (�	      �   ,�	      �   0�	      �   4�	      �   8�	        <�	      %  @�	      M  D�	      ~  H�	      �  P�	      �  T�	      �  X�	      �  \�	      �  `�	        d�	      B  h�	      Z  l�	      q  p�	      �  t�	      �  x�	      �  |�	      �  ��	      
  ��	      5  ��	      d  ��	      �  ��	      �  ��	      �  ��	      �  ��	      �  ��	      �  ��	        ��	        ��	      "  ��	      0  ��	      D  ��	      X  ��	      o  ��	      }  ��	      �  ��	      �  ��	      �  ��	      �  ��	      �  ��	      �  ��	      �  ��	        ��	        ��	      +  ��	      @  ��	      U  ��	      i  ��	      x  ��	      �   �	      �  �	      �  �	      �  �	      �  �	      �  �	        �	      1  �	      Q   �	      m  $�	      �  (�	      �  ,�	      �  0�	      �  4�	        8�	        <�	      <  @�	      R  D�	      j  H�	      �  L�	      �  P�	      �  T�	      �  X�	      �  \�	        `�	      9  d�	      X  h�	      w  l�	      �  p�	      �  t�	      �  x�	      �  |�	      	  ��	      E	  ��	      p	  ��	      �	  ��	      �	  ��	      z
  ,D      �
        �
  8D     
 �
  ��      �
           ���
           ���
  �@     �
  0�K       ��    =  ���     f   �s     �  ��p     �  �               ��           ��(   �P     n           ��y           ���           ���           ���           ���  ��2     �  ��@     �  ���                ��'           ��0           ��<  ���    [           ��g           ��t           ���  ��"     �           ���  �E     �           ���           ���  �E     2           ��D           ��P           ��[           ��o           ��           ���  Ќ2     �           ���  0�$     �           ���           ��           ��           ��'           ��2           ��@  F     P           ��\           ��l           ��u           ���           ���           ���           ���           ���  �G     �  �G     �  F     �  @F@               ��           ��(           ��7           ��?           ��J           ��\           ��r           ���  �O     �           ���           ���           ���   �(       �U     O   U8     l  `U8     �  �U     �  �U     �   S     �  �R     �  �R        Rh     ;  �R     X  �R     u  �R     �   QD     �  �R     �  �QD       �R     &  �R     F  �R     f   P�     �  �R     �  �R     �  xR     �  hR     	  �U     +  `�'     P  �U     l           ��{           ���           ���           ���           ���           ���           ���           ���  S       �	�                 ��4           ��A           ��N  �	     n           ��~           ���           ���           ���  �#     �  �#       � 	$     1  �#     ^  �#!     �  �%    �  [     �  �D     1  @ 	)     ]  l 	     �           ���  @'     �  P'     �  �'     )  �'     V  �'     �  �'     �  �'     �  �'       �')     A   ()     v  �D     �  �D     �  ��2     �   !	*     )  @!	)     U  l!	     �  x!	     �  �!	$     �   "	$                ��  [     8           ��I           ��W  �)�     c  �*F     o  �*      �+[     �  P,�    �   -	�     �   .h     �  �.o     �   /t     �  �/S     �  �/?        0U       �0#     (  �0�     6  �1}     D  2q     f  �2i     r   3�     �  �3�     �  �4�     �  @5�'    �  �o�     �  pp2    �   2	�    �  �\.      �g�    #  `j&    A  �m5    V   d�    g  �q`    v   �4    }  ��$    �  s�    �  ��    �  ��    �  ���    �  ��7    �   �#    �  ��[     �  ���    �  `��       @�d        .	�    3  �D    T           ��T           ��^           ��k  ��A     x   ��	    �   ��    �  � �    �  [     �  ��    �  PD    �  �t     �   �       ��     7  ��    L       ^  ��       c  ��       h  ��       n  �       t  �	       z  ��         b�       �  ��       �  ��       �  ��       �  B�       �  ��       �  ��       �  �       �  {�       �  ��       �  ��       �  C�       �  ��       �  ��       �  �       �  r�       �  ��       �  .�       �  Q�       �  ��       �  *�       �  ��       �  ��       �  �       �  e�       �  \�          H�          ��          ��          @�          ��          ��       "   {�       (   ��       .   ��       4   ��       :   Z�       @   ��       F   Q�       L   ��       R   ��       X   0       ^           d          j           p   �       v   �       |   p       �   0       �          �   �       �   �       �   �       �   �       �   �       �   �       �   `       �   0       �           �   �       �   �       �   p       �           �   `       �   �       �   p       �          �   <       �   0        !  �       !         !  $       !  �       !  �       !  �       $!  �       *!  ?       0!  I       6!  R       <!  [       B!  d       H!  m       N!  v       T!         Z!  �       `!  �       f!  �       l!  �       r!  �       x!  @       ~!         �!  @
       �!  �	       �!  �
       �!           ��k  �A     �!  �     �!  ��     �!  ��     �!  `w     �!  �h     "  P/    "  �{     ;"       L"  f    f"  �'    o"  � I    �"   "�     �"  �"n    �"  4[     �"  0[     �"  @[     �"  <[     �"  P       �"  �       �"         �"  @       �"  �       �"  �       #  �       #           ��2#  �       7#           ��F#  ��     a#  4�
     |#  <E     �#  :�A     �#  k�     �#  l�     �#  m�     �#  n�     $  o�     2$  p�     C$  t�     T$  x�     e$  |�     |$  ��     �$  ��     �$  ��     �$  ��     �$  ��     �$  ��     %  ��     L%  ��     �%  ��     �%  ��     �%  ��     �%  ��     �%  ��     &  ��     =&  ��     i&  ��     �&  ��     �&  ��     �&  ��     �&  ��     �&  ��     )'  ��     T'  ��     �'  ��     �'  ��     �'  ��     (  ��     %(  ��     <(  ��     O(  ��     a(  ��     y(   �     �(  �     �(  �     �(  �     �(  �     �(  �     )  �     )  �     +)   �     D)  $�     ])  (�     p)  ,�     �)  0�     �)  4�     �)  8�     �)  <�     �)  @�     �)  D�     *  H�     +*  L�     D*  P�     X*  T�     m*  X�     �*  \�     �*  `�     �*  d�     �*  h�     �*  l�     +  p�     9+  t�     ^+  x�     +  |�     �+  ��     �+  ��     �+  ��     ,  ��     2,  ��     O,  ��     q,  ��     �,  ��     �,  ��     �,  ��     �,  ��     -  ��     --  ��     Q-  ��     t-  ��     �-  ��     �-  ��     �-  ��     .  ��     ,.  ��     S.  ��     {.  ��     �.  ��     �.  ��     �.  ��     '/  ��     G/  ��     g/  {�     �/           ��F#  ��     a#  ��
     |#  =E     �#  ��A     �#  
�     �#  �     �#  �     �#  �     $  �     2$  �     C$  �     T$  �     e$  �     |$   �     �$  $�     �$  (�     �$  ,�     �$  0�     �$  4�     %  8�     L%  <�     �%  @�     �%  H�     �%  L�     �%  P�     �%  T�     &  X�     =&  \�     i&  `�     �&  d�     �&  h�     �&  l�     �&  p�     �&  t�     )'  x�     T'  |�     �'  ��     �'  ��     �'  ��     (  ��     %(  ��     <(  ��     O(  ��     a(  ��     y(  ��     �(  ��     �(  ��     �(  ��     �(  ��     �(  ��     )  ��     )  ��     +)  ��     D)  ��     ])  ��     p)  ��     �)  ��     �)  ��     �)  ��     �)  ��     �)  ��     �)  ��     *  ��     +*  ��     D*  ��     X*  ��     m*  ��     �*  ��     �*   �     �*  �     �*  �     �*  �     +  �     9+  �     ^+  �     +  �     �+   �     �+  $�     �+  (�     ,  ,�     2,  0�     O,  4�     q,  8�     �,  <�     �,  @�     �,  D�     �,  H�     -  L�     --  P�     Q-  T�     t-  X�     �-  \�     �-  `�     �-  d�     .  h�     ,.  l�     S.  p�     {.  t�     �.  x�     �.  |�     �.  ��     '/  ��     G/  ��     �/  9�     �/           ��F#  ��     a#  S�
     |#  >E     �#  ]�A     �#  ��     �#  ��     �#  ��     �#  ��     $  ��     2$  ��     C$  ��     T$  ��     e$  ��     |$  ��     �$  ��     �$  ��     �$  ��     �$  ��     �$  ��     %  ��     L%  ��     �%  ��     �%  ��     �%  ��     �%  ��     �%  ��     &  ��     =&  ��     i&  ��     �&  ��     �&  ��     �&  ��     �&  ��     �&  ��     )'   �     T'  �     �'  �     �'  �     �'  �     (  �     %(  �     <(  �     O(   �     a(  $�     y(  (�     �(  ,�     �(  0�     �(  4�     �(  8�     �(  <�     )  @�     )  D�     +)  H�     D)  L�     ])  P�     p)  T�     �)  X�     �)  \�     �)  `�     �)  d�     �)  h�     �)  l�     *  p�     +*  t�     D*  x�     X*  |�     m*  ��     �*  ��     �*  ��     �*  ��     �*  ��     �*  ��     +  ��     9+  ��     ^+  ��     +  ��     �+  ��     �+  ��     �+  ��     ,  ��     2,  ��     O,  ��     q,  ��     �,  ��     �,  ��     �,  ��     �,  ��     -  ��     --  ��     Q-  ��     t-  ��     �-  ��     �-  ��     �-  ��     .  ��     ,.  ��     S.  ��     {.  ��     �.   �     �.  �     �.  �     '/  �     G/  �     �/  ��     0           ��F#  �     a#  ��
     |#  ?E     �#  ��A     �#  1�     �#  2�     �#  3�     �#  4�     $  5�     2$  8�     C$  <�     T$  @�     e$  D�     |$  H�     �$  L�     �$  P�     �$  T�     �$  X�     �$  \�     %  `�     L%  d�     �%  h�     �%  p�     �%  t�     �%  x�     �%  |�     &  ��     =&  ��     i&  ��     �&  ��     �&  ��     �&  ��     �&  ��     �&  ��     )'  ��     T'  ��     �'  ��     �'  ��     �'  ��     (  ��     %(  ��     <(  ��     O(  ��     a(  ��     y(  ��     �(  ��     �(  ��     �(  ��     �(  ��     �(  ��     )  ��     )  ��     +)  ��     D)  ��     ])  ��     p)  ��     �)  ��     �)  ��     �)   �     �)  �     �)  �     �)  �     *  �     +*  �     D*  �     X*  �     m*   �     �*  $�     �*  (�     �*  ,�     �*  0�     �*  4�     +  8�     9+  <�     ^+  @�     +  D�     �+  H�     �+  L�     �+  P�     ,  T�     2,  X�     O,  \�     q,  `�     �,  d�     �,  h�     �,  l�     �,  p�     -  t�     --  x�     Q-  |�     t-  ��     �-  ��     �-  ��     �-  ��     .  ��     ,.  ��     S.  ��     {.  ��     �.  ��     �.  ��     �.  ��     '/  ��     G/  ��     0  6�     80           ��F#  ��     a#  P�
     �#  ��     �#  ��     �#  ��     �#  ��     $  ��     2$  ��     C$  ��     T$  ��     e$  ��     |$  ��     �$  ��     �$  ��     �$  ��     �$  ��     �$  ��     %  ��     L%  ��     �%  ��     �%  ��     �%  ��     �%   �     �%  �     &  �     =&  �     i&  �     �&  �     �&  �     �&  �     �&   �     �&  $�     )'  (�     T'  ,�     �'  0�     �'  4�     �'  8�     (  <�     %(  @�     <(  D�     O(  H�     a(  L�     y(  P�     �(  T�     �(  X�     �(  \�     �(  `�     �(  d�     )  h�     )  l�     +)  p�     D)  t�     ])  x�     p)  |�     �)  ��     �)  ��     �)  ��     �)  ��     �)  ��     �)  ��     *  ��     +*  ��     D*  ��     X*  ��     m*  ��     �*  ��     �*  ��     �*  ��     �*  ��     �*  ��     +  ��     9+  ��     ^+  ��     +  ��     �+  ��     �+  ��     �+  ��     ,  ��     2,  ��     O,  ��     q,  ��     �,  ��     �,  ��     �,  ��     �,  ��     -  ��     --   �     Q-  �     t-  �     �-  �     �-  �     �-  �     .  �     ,.  �     S.   �     {.  $�     �.  (�     �.  ,�     �.  0�     '/  4�     G/  8�     C0           ��F#  @�     a#  �
     2$  D�     C$  H�     T$  L�     e$  P�     |$  T�     �$  X�     �$  \�     �$  `�     �$  d�     �$  h�     %  l�     L%  p�     �%  x�     �%  ��     �%  ��     �%  ��     �%  ��     &  ��     =&  ��     i&  ��     �&  ��     �&  ��     �&  ��     �&  ��     �&  ��     )'  ��     T'  ��     �'  ��     �'  ��     �'  ��     (  ��     %(  ��     <(  ��     O(  ��     a(  ��     y(  ��     �(  ��     �(  ��     �(  ��     �(  ��     �(  ��     )  ��     )  ��     +)  ��     D)  ��     ])   �     p)  �     �)  �     �)  �     �)  �     �)  �     �)  �     �)  �     *   �     +*  $�     D*  (�     X*  ,�     m*  0�     �*  4�     �*  8�     �*  <�     �*  @�     �*  D�     +  H�     9+  L�     ^+  P�     +  T�     �+  X�     �+  \�     �+  `�     ,  d�     2,  h�     O,  l�     q,  p�     �,  t�     �,  x�     �,  |�     �,  ��     �#  ��     �#  ��     �#  ��     �#  ��     $  ��     -  ��     --  ��     Q-  ��     t-  ��     �-  ��     �-  ��     �-  ��     .  ��     ,.  ��     S.  ��     {.  ��     �.  ��     �.  ��     �.  ��     '/  ��     G/  ��     M0           ��`0           ��s0           ���0           ���#  �@	     �#  �@	     �#  �@	     �#  �@	     $  �@	     2$  �@	     C$  �@	     T$  �@	     e$  �@	     |$  �@	     �$  �@	     �$  �@	     �$  �@	     �$  �@	     �$  �@	     %  �@	     L%  �@	     �%  �@	     �%  �@	     �%  �@	     �%   A	     �%  A	     &  A	     =&  A	     i&  A	     �&  A	     �&  A	     �&  A	     �&   A	     �&  $A	     )'  (A	     T'  ,A	     �'  0A	     �'  4A	     �'  8A	     (  <A	     %(  @A	     <(  DA	     O(  HA	     a(  LA	     y(  PA	     �(  TA	     �(  XA	     �(  \A	     �(  `A	     �(  dA	     )  hA	     )  lA	     +)  pA	     D)  tA	     ])  xA	     p)  |A	     �)  �A	     �)  �A	     �)  �A	     �)  �A	     �)  �A	     �)  �A	     *  �A	     +*  �A	     D*  �A	     X*  �A	     m*  �A	     �*  �A	     �*  �A	     �*  �A	     �*  �A	     �*  �A	     +  �A	     9+  �A	     ^+  �A	     +  �A	     �+  �A	     �+  �A	     �+  �A	     ,  �A	     2,  �A	     O,  �A	     q,  �A	     �,  �A	     �,  �A	     �,  �A	     �,  �A	     -  �A	     --   B	     Q-  B	     t-  B	     �-  B	     �-  B	     �-  B	     .  B	     ,.  B	     S.   B	     {.  $B	     �.  (B	     �.  ,B	     �.  0B	     '/  4B	     G/  8B	     �0           ���#  @B	     �#  AB	     �#  BB	     �#  CB	     $  DB	     2$  HB	     C$  LB	     T$  PB	     e$  TB	     |$  XB	     �$  \B	     �$  `B	     �$  dB	     �$  hB	     �$  lB	     %  pB	     L%  tB	     �%  xB	     �%  �B	     �%  �B	     �%  �B	     �%  �B	     &  �B	     =&  �B	     i&  �B	     �&  �B	     �&  �B	     �&  �B	     �&  �B	     �&  �B	     )'  �B	     T'  �B	     �'  �B	     �'  �B	     �'  �B	     (  �B	     %(  �B	     <(  �B	     O(  �B	     a(  �B	     y(  �B	     �(  �B	     �(  �B	     �(  �B	     �(  �B	     �(  �B	     )  �B	     )  �B	     +)  �B	     D)  �B	     ])   C	     p)  C	     �)  C	     �)  C	     �)  C	     �)  C	     �)  C	     �)  C	     *   C	     +*  $C	     D*  (C	     X*  ,C	     m*  0C	     �*  4C	     �*  8C	     �*  <C	     �*  @C	     �*  DC	     +  HC	     9+  LC	     ^+  PC	     +  TC	     �+  XC	     �+  \C	     �+  `C	     ,  dC	     2,  hC	     O,  lC	     q,  pC	     �,  tC	     �,  xC	     �,  |C	     �,  �C	     -  �C	     --  �C	     Q-  �C	     t-  �C	     �-  �C	     �-  �C	     �-  �C	     .  �C	     ,.  �C	     S.  �C	     {.  �C	     �.  �C	     �.  �C	     �.  �C	     '/  �C	     G/  �C	     �0           ���#  �C	     �#  �C	     �#  �C	     �#  �C	     $  �C	     2$  �C	     C$  �C	     T$  �C	     e$  �C	     |$  �C	     �$  �C	     �$  �C	     �$  �C	     �$  �C	     �$  �C	     %  �C	     L%  �C	     �%   D	     �%  D	     �%  D	     �%  D	     �%  D	     &  D	     =&  D	     i&   D	     �&  $D	     �&  (D	     �&  ,D	     �&  0D	     �&  4D	     )'  8D	     T'  <D	     �'  @D	     �'  DD	     �'  HD	     (  LD	     %(  PD	     <(  TD	     O(  XD	     a(  \D	     y(  `D	     �(  dD	     �(  hD	     �(  lD	     �(  pD	     �(  tD	     )  xD	     )  |D	     +)  �D	     D)  �D	     ])  �D	     p)  �D	     �)  �D	     �)  �D	     �)  �D	     �)  �D	     �)  �D	     �)  �D	     *  �D	     +*  �D	     D*  �D	     X*  �D	     m*  �D	     �*  �D	     �*  �D	     �*  �D	     �*  �D	     �*  �D	     +  �D	     9+  �D	     ^+  �D	     +  �D	     �+  �D	     �+  �D	     �+  �D	     ,  �D	     2,  �D	     O,  �D	     q,  �D	     �,  �D	     �,   E	     �,  E	     �,  E	     -  E	     --  E	     Q-  E	     t-  E	     �-  E	     �-   E	     �-  $E	     .  (E	     ,.  ,E	     S.  0E	     {.  4E	     �.  8E	     �.  <E	     �.  @E	     '/  DE	     G/  HE	     �0           ���#  PE	     �#  QE	     �#  RE	     �#  SE	     $  TE	     2$  XE	     C$  \E	     T$  `E	     e$  dE	     |$  hE	     �$  lE	     �$  pE	     �$  tE	     �$  xE	     �$  |E	     %  �E	     L%  �E	     �%  �E	     �%  �E	     �%  �E	     �%  �E	     �%  �E	     &  �E	     =&  �E	     i&  �E	     �&  �E	     �&  �E	     �&  �E	     �&  �E	     �&  �E	     )'  �E	     T'  �E	     �'  �E	     �'  �E	     �'  �E	     (  �E	     %(  �E	     <(  �E	     O(  �E	     a(  �E	     y(  �E	     �(  �E	     �(  �E	     �(  �E	     �(  �E	     �(  �E	     )   F	     )  F	     +)  F	     D)  F	     ])  F	     p)  F	     �)  F	     �)  F	     �)   F	     �)  $F	     �)  (F	     �)  ,F	     *  0F	     +*  4F	     D*  8F	     X*  <F	     m*  @F	     �*  DF	     �*  HF	     �*  LF	     �*  PF	     �*  TF	     +  XF	     9+  \F	     ^+  `F	     +  dF	     �+  hF	     �+  lF	     �+  pF	     ,  tF	     2,  xF	     O,  |F	     q,  �F	     �,  �F	     �,  �F	     �,  �F	     �,  �F	     -  �F	     --  �F	     Q-  �F	     t-  �F	     �-  �F	     �-  �F	     �-  �F	     .  �F	     ,.  �F	     S.  �F	     {.  �F	     �.  �F	     �.  �F	     �.  �F	     '/  �F	     G/  �F	     �0           ���#  �F	     �#  �F	     �#  �F	     �#  �F	     $  �F	     2$  �F	     C$  �F	     T$  �F	     e$  �F	     |$  �F	     �$  �F	     �$  �F	     �$  �F	     �$   G	     �$  G	     %  G	     L%  G	     �%  G	     �%  G	     �%  G	     �%   G	     �%  $G	     &  (G	     =&  ,G	     i&  0G	     �&  4G	     �&  8G	     �&  <G	     �&  @G	     �&  DG	     )'  HG	     T'  LG	     �'  PG	     �'  TG	     �'  XG	     (  \G	     %(  `G	     <(  dG	     O(  hG	     a(  lG	     y(  pG	     �(  tG	     �(  xG	     �(  |G	     �(  �G	     �(  �G	     )  �G	     )  �G	     +)  �G	     D)  �G	     ])  �G	     p)  �G	     �)  �G	     �)  �G	     �)  �G	     �)  �G	     �)  �G	     �)  �G	     *  �G	     +*  �G	     D*  �G	     X*  �G	     m*  �G	     �*  �G	     �*  �G	     �*  �G	     �*  �G	     �*  �G	     +  �G	     9+  �G	     ^+  �G	     +  �G	     �+  �G	     �+  �G	     �+  �G	     ,  �G	     2,   H	     O,  H	     q,  H	     �,  H	     �,  H	     �,  H	     �,  H	     -  H	     --   H	     Q-  $H	     t-  (H	     �-  ,H	     �-  0H	     �-  4H	     .  8H	     ,.  <H	     S.  @H	     {.  DH	     �.  HH	     �.  LH	     �.  PH	     '/  TH	     G/  XH	     �0           ���#  `H	     �#  aH	     �#  bH	     �#  cH	     $  dH	     2$  hH	     C$  lH	     T$  pH	     e$  tH	     |$  xH	     �$  |H	     �$  �H	     �$  �H	     �$  �H	     �$  �H	     %  �H	     L%  �H	     �%  �H	     �%  �H	     �%  �H	     �%  �H	     �%  �H	     &  �H	     =&  �H	     i&  �H	     �&  �H	     �&  �H	     �&  �H	     �&  �H	     �&  �H	     )'  �H	     T'  �H	     �'  �H	     �'  �H	     �'  �H	     (  �H	     %(  �H	     <(  �H	     O(  �H	     a(  �H	     y(  �H	     �(  �H	     �(   I	     �(  I	     �(  I	     �(  I	     )  I	     )  I	     +)  I	     D)  I	     ])   I	     p)  $I	     �)  (I	     �)  ,I	     �)  0I	     �)  4I	     �)  8I	     �)  <I	     *  @I	     +*  DI	     D*  HI	     X*  LI	     m*  PI	     �*  TI	     �*  XI	     �*  \I	     �*  `I	     �*  dI	     +  hI	     9+  lI	     ^+  pI	     +  tI	     �+  xI	     �+  |I	     �+  �I	     ,  �I	     2,  �I	     O,  �I	     q,  �I	     �,  �I	     �,  �I	     �,  �I	     �,  �I	     -  �I	     --  �I	     Q-  �I	     t-  �I	     �-  �I	     �-  �I	     �-  �I	     .  �I	     ,.  �I	     S.  �I	     {.  �I	     �.  �I	     �.  �I	     �.  �I	     '/  �I	     G/  �I	     �0           ���#  �I	     �#  �I	     �#  �I	     �#  �I	     $  �I	     2$  �I	     C$  �I	     T$  �I	     e$  �I	     |$   J	     �$  J	     �$  J	     �$  J	     �$  J	     �$  J	     %  J	     L%  J	     �%   J	     �%  (J	     �%  ,J	     �%  0J	     �%  4J	     &  8J	     =&  <J	     i&  @J	     �&  DJ	     �&  HJ	     �&  LJ	     �&  PJ	     �&  TJ	     )'  XJ	     T'  \J	     �'  `J	     �'  dJ	     �'  hJ	     (  lJ	     %(  pJ	     <(  tJ	     O(  xJ	     a(  |J	     y(  �J	     �(  �J	     �(  �J	     �(  �J	     �(  �J	     �(  �J	     )  �J	     )  �J	     +)  �J	     D)  �J	     ])  �J	     p)  �J	     �)  �J	     �)  �J	     �)  �J	     �)  �J	     �)  �J	     �)  �J	     *  �J	     +*  �J	     D*  �J	     X*  �J	     m*  �J	     �*  �J	     �*  �J	     �*  �J	     �*  �J	     �*  �J	     +  �J	     9+  �J	     ^+  �J	     +  �J	     �+   K	     �+  K	     �+  K	     ,  K	     2,  K	     O,  K	     q,  K	     �,  K	     �,   K	     �,  $K	     �,  (K	     -  ,K	     --  0K	     Q-  4K	     t-  8K	     �-  <K	     �-  @K	     �-  DK	     .  HK	     ,.  LK	     S.  PK	     {.  TK	     �.  XK	     �.  \K	     �.  `K	     '/  dK	     G/  hK	     �0           ���#  pK	     �#  qK	     �#  rK	     �#  sK	     $  tK	     2$  xK	     C$  |K	     T$  �K	     e$  �K	     |$  �K	     �$  �K	     �$  �K	     �$  �K	     �$  �K	     �$  �K	     %  �K	     L%  �K	     �%  �K	     �%  �K	     �%  �K	     �%  �K	     �%  �K	     &  �K	     =&  �K	     i&  �K	     �&  �K	     �&  �K	     �&  �K	     �&  �K	     �&  �K	     )'  �K	     T'  �K	     �'  �K	     �'  �K	     �'  �K	     (  �K	     %(  �K	     <(  �K	     O(   L	     a(  L	     y(  L	     �(  L	     �(  L	     �(  L	     �(  L	     �(  L	     )   L	     )  $L	     +)  (L	     D)  ,L	     ])  0L	     p)  4L	     �)  8L	     �)  <L	     �)  @L	     �)  DL	     �)  HL	     �)  LL	     *  PL	     +*  TL	     D*  XL	     X*  \L	     m*  `L	     �*  dL	     �*  hL	     �*  lL	     �*  pL	     �*  tL	     +  xL	     9+  |L	     ^+  �L	     +  �L	     �+  �L	     �+  �L	     �+  �L	     ,  �L	     2,  �L	     O,  �L	     q,  �L	     �,  �L	     �,  �L	     �,  �L	     �,  �L	     -  �L	     --  �L	     Q-  �L	     t-  �L	     �-  �L	     �-  �L	     �-  �L	     .  �L	     ,.  �L	     S.  �L	     {.  �L	     �.  �L	     �.  �L	     �.  �L	     '/  �L	     G/  �L	     1           ���#  �L	     �#  �L	     �#  �L	     �#  �L	     $  �L	     2$   M	     C$  M	     T$  M	     e$  M	     |$  M	     �$  M	     �$  M	     �$  M	     �$   M	     �$  $M	     %  (M	     L%  ,M	     �%  0M	     �%  8M	     �%  <M	     �%  @M	     �%  DM	     &  HM	     =&  LM	     i&  PM	     �&  TM	     �&  XM	     �&  \M	     �&  `M	     �&  dM	     )'  hM	     T'  lM	     �'  pM	     �'  tM	     �'  xM	     (  |M	     %(  �M	     <(  �M	     O(  �M	     a(  �M	     y(  �M	     �(  �M	     �(  �M	     �(  �M	     �(  �M	     �(  �M	     )  �M	     )  �M	     +)  �M	     D)  �M	     ])  �M	     p)  �M	     �)  �M	     �)  �M	     �)  �M	     �)  �M	     �)  �M	     �)  �M	     *  �M	     +*  �M	     D*  �M	     X*  �M	     m*  �M	     �*  �M	     �*  �M	     �*  �M	     �*  �M	     �*  �M	     +   N	     9+  N	     ^+  N	     +  N	     �+  N	     �+  N	     �+  N	     ,  N	     2,   N	     O,  $N	     q,  (N	     �,  ,N	     �,  0N	     �,  4N	     �,  8N	     -  <N	     --  @N	     Q-  DN	     t-  HN	     �-  LN	     �-  PN	     �-  TN	     .  XN	     ,.  \N	     S.  `N	     {.  dN	     �.  hN	     �.  lN	     �.  pN	     '/  tN	     G/  xN	      1           ���#  �N	     �#  �N	     �#  �N	     �#  �N	     $  �N	     2$  �N	     C$  �N	     T$  �N	     e$  �N	     |$  �N	     �$  �N	     �$  �N	     �$  �N	     �$  �N	     �$  �N	     %  �N	     L%  �N	     �%  �N	     �%  �N	     �%  �N	     �%  �N	     �%  �N	     &  �N	     =&  �N	     i&  �N	     �&  �N	     �&  �N	     �&  �N	     �&  �N	     �&  �N	     )'  �N	     T'  �N	     �'  �N	     �'  �N	     �'   O	     (  O	     %(  O	     <(  O	     O(  O	     a(  O	     y(  O	     �(  O	     �(   O	     �(  $O	     �(  (O	     �(  ,O	     )  0O	     )  4O	     +)  8O	     D)  <O	     ])  @O	     p)  DO	     �)  HO	     �)  LO	     �)  PO	     �)  TO	     �)  XO	     �)  \O	     *  `O	     +*  dO	     D*  hO	     X*  lO	     m*  pO	     �*  tO	     �*  xO	     �*  |O	     �*  �O	     �*  �O	     +  �O	     9+  �O	     ^+  �O	     +  �O	     �+  �O	     �+  �O	     �+  �O	     ,  �O	     2,  �O	     O,  �O	     q,  �O	     �,  �O	     �,  �O	     �,  �O	     �,  �O	     -  �O	     --  �O	     Q-  �O	     t-  �O	     �-  �O	     �-  �O	     �-  �O	     .  �O	     ,.  �O	     S.  �O	     {.  �O	     �.  �O	     �.  �O	     �.  �O	     '/  �O	     G/   P	     01           ���#  P	     �#  	P	     �#  
P	     �#  P	     $  P	     2$  P	     C$  P	     T$  P	     e$  P	     |$   P	     �$  $P	     �$  (P	     �$  ,P	     �$  0P	     �$  4P	     %  8P	     L%  <P	     �%  @P	     �%  HP	     �%  LP	     �%  PP	     �%  TP	     &  XP	     =&  \P	     i&  `P	     �&  dP	     �&  hP	     �&  lP	     �&  pP	     �&  tP	     )'  xP	     T'  |P	     �'  �P	     �'  �P	     �'  �P	     (  �P	     %(  �P	     <(  �P	     O(  �P	     a(  �P	     y(  �P	     �(  �P	     �(  �P	     �(  �P	     �(  �P	     �(  �P	     )  �P	     )  �P	     +)  �P	     D)  �P	     ])  �P	     p)  �P	     �)  �P	     �)  �P	     �)  �P	     �)  �P	     �)  �P	     �)  �P	     *  �P	     +*  �P	     D*  �P	     X*  �P	     m*  �P	     �*  �P	     �*   Q	     �*  Q	     �*  Q	     �*  Q	     +  Q	     9+  Q	     ^+  Q	     +  Q	     �+   Q	     �+  $Q	     �+  (Q	     ,  ,Q	     2,  0Q	     O,  4Q	     q,  8Q	     �,  <Q	     �,  @Q	     �,  DQ	     �,  HQ	     -  LQ	     --  PQ	     Q-  TQ	     t-  XQ	     �-  \Q	     �-  `Q	     �-  dQ	     .  hQ	     ,.  lQ	     S.  pQ	     {.  tQ	     �.  xQ	     �.  |Q	     �.  �Q	     '/  �Q	     G/  �Q	     H1           ���#  �Q	     �#  �Q	     �#  �Q	     �#  �Q	     $  �Q	     2$  �Q	     C$  �Q	     T$  �Q	     e$  �Q	     |$  �Q	     �$  �Q	     �$  �Q	     �$  �Q	     �$  �Q	     �$  �Q	     %  �Q	     L%  �Q	     �%  �Q	     �%  �Q	     �%  �Q	     �%  �Q	     �%  �Q	     &  �Q	     =&  �Q	     i&  �Q	     �&  �Q	     �&  �Q	     �&  �Q	     �&  �Q	     �&  �Q	     )'   R	     T'  R	     �'  R	     �'  R	     �'  R	     (  R	     %(  R	     <(  R	     O(   R	     a(  $R	     y(  (R	     �(  ,R	     �(  0R	     �(  4R	     �(  8R	     �(  <R	     )  @R	     )  DR	     +)  HR	     D)  LR	     ])  PR	     p)  TR	     �)  XR	     �)  \R	     �)  `R	     �)  dR	     �)  hR	     �)  lR	     *  pR	     +*  tR	     D*  xR	     X*  |R	     m*  �R	     �*  �R	     �*  �R	     �*  �R	     �*  �R	     �*  �R	     +  �R	     9+  �R	     ^+  �R	     +  �R	     �+  �R	     �+  �R	     �+  �R	     ,  �R	     2,  �R	     O,  �R	     q,  �R	     �,  �R	     �,  �R	     �,  �R	     �,  �R	     -  �R	     --  �R	     Q-  �R	     t-  �R	     �-  �R	     �-  �R	     �-  �R	     .  �R	     ,.  �R	     S.  �R	     {.  �R	     �.   S	     �.  S	     �.  S	     '/  S	     G/  S	     U1           ���#  S	     �#  S	     �#  S	     �#  S	     $  S	     2$   S	     C$  $S	     T$  (S	     e$  ,S	     |$  0S	     �$  4S	     �$  8S	     �$  <S	     �$  @S	     �$  DS	     %  HS	     L%  LS	     �%  PS	     �%  XS	     �%  \S	     �%  `S	     �%  dS	     &  hS	     =&  lS	     i&  pS	     �&  tS	     �&  xS	     �&  |S	     �&  �S	     �&  �S	     )'  �S	     T'  �S	     �'  �S	     �'  �S	     �'  �S	     (  �S	     %(  �S	     <(  �S	     O(  �S	     a(  �S	     y(  �S	     �(  �S	     �(  �S	     �(  �S	     �(  �S	     �(  �S	     )  �S	     )  �S	     +)  �S	     D)  �S	     ])  �S	     p)  �S	     �)  �S	     �)  �S	     �)  �S	     �)  �S	     �)  �S	     �)  �S	     *  �S	     +*  �S	     D*   T	     X*  T	     m*  T	     �*  T	     �*  T	     �*  T	     �*  T	     �*  T	     +   T	     9+  $T	     ^+  (T	     +  ,T	     �+  0T	     �+  4T	     �+  8T	     ,  <T	     2,  @T	     O,  DT	     q,  HT	     �,  LT	     �,  PT	     �,  TT	     �,  XT	     -  \T	     --  `T	     Q-  dT	     t-  hT	     �-  lT	     �-  pT	     �-  tT	     .  xT	     ,.  |T	     S.  �T	     {.  �T	     �.  �T	     �.  �T	     �.  �T	     '/  �T	     G/  �T	     a1           ���#  �T	     �#  �T	     �#  �T	     �#  �T	     $  �T	     2$  �T	     C$  �T	     T$  �T	     e$  �T	     |$  �T	     �$  �T	     �$  �T	     �$  �T	     �$  �T	     �$  �T	     %  �T	     L%  �T	     �%  �T	     �%  �T	     �%  �T	     �%  �T	     �%  �T	     &  �T	     =&  �T	     i&  �T	     �&  �T	     �&   U	     �&  U	     �&  U	     �&  U	     )'  U	     T'  U	     �'  U	     �'  U	     �'   U	     (  $U	     %(  (U	     <(  ,U	     O(  0U	     a(  4U	     y(  8U	     �(  <U	     �(  @U	     �(  DU	     �(  HU	     �(  LU	     )  PU	     )  TU	     +)  XU	     D)  \U	     ])  `U	     p)  dU	     �)  hU	     �)  lU	     �)  pU	     �)  tU	     �)  xU	     �)  |U	     *  �U	     +*  �U	     D*  �U	     X*  �U	     m*  �U	     �*  �U	     �*  �U	     �*  �U	     �*  �U	     �*  �U	     +  �U	     9+  �U	     ^+  �U	     +  �U	     �+  �U	     �+  �U	     �+  �U	     ,  �U	     2,  �U	     O,  �U	     q,  �U	     �,  �U	     �,  �U	     �,  �U	     �,  �U	     -  �U	     --  �U	     Q-  �U	     t-  �U	     �-  �U	     �-  �U	     �-  �U	     .   V	     ,.  V	     S.  V	     {.  V	     �.  V	     �.  V	     �.  V	     '/  V	     G/   V	     t1           ���#  (V	     �#  )V	     �#  *V	     �#  +V	     $  ,V	     2$  0V	     C$  4V	     T$  8V	     e$  <V	     |$  @V	     �$  DV	     �$  HV	     �$  LV	     �$  PV	     �$  TV	     %  XV	     L%  \V	     �%  `V	     �%  hV	     �%  lV	     �%  pV	     �%  tV	     &  xV	     =&  |V	     i&  �V	     �&  �V	     �&  �V	     �&  �V	     �&  �V	     �&  �V	     )'  �V	     T'  �V	     �'  �V	     �'  �V	     �'  �V	     (  �V	     %(  �V	     <(  �V	     O(  �V	     a(  �V	     y(  �V	     �(  �V	     �(  �V	     �(  �V	     �(  �V	     �(  �V	     )  �V	     )  �V	     +)  �V	     D)  �V	     ])  �V	     p)  �V	     �)  �V	     �)  �V	     �)  �V	     �)  �V	     �)   W	     �)  W	     *  W	     +*  W	     D*  W	     X*  W	     m*  W	     �*  W	     �*   W	     �*  $W	     �*  (W	     �*  ,W	     +  0W	     9+  4W	     ^+  8W	     +  <W	     �+  @W	     �+  DW	     �+  HW	     ,  LW	     2,  PW	     O,  TW	     q,  XW	     �,  \W	     �,  `W	     �,  dW	     �,  hW	     -  lW	     --  pW	     Q-  tW	     t-  xW	     �-  |W	     �-  �W	     �-  �W	     .  �W	     ,.  �W	     S.  �W	     {.  �W	     �.  �W	     �.  �W	     �.  �W	     '/  �W	     G/  �W	     �1           ���1           ���1           ���1           ���1           ���1           ���1           ���1           ���1           ���1           ���1           ��
2           ��2           �� 2           ��<2           ��J2           ���#  �W	     �#  �W	     �#  �W	     �#  �W	     $  �W	     2$  �W	     C$  �W	     T$  �W	     e$  �W	     |$  �W	     �$  �W	     �$  �W	     �$  �W	     �$   X	     �$  X	     %  X	     L%  X	     �%  X	     �%  X	     �%  X	     �%   X	     �%  $X	     &  (X	     =&  ,X	     i&  0X	     �&  4X	     �&  8X	     �&  <X	     �&  @X	     �&  DX	     )'  HX	     T'  LX	     �'  PX	     �'  TX	     �'  XX	     (  \X	     %(  `X	     <(  dX	     O(  hX	     a(  lX	     y(  pX	     �(  tX	     �(  xX	     �(  |X	     �(  �X	     �(  �X	     )  �X	     )  �X	     +)  �X	     D)  �X	     ])  �X	     p)  �X	     �)  �X	     �)  �X	     �)  �X	     �)  �X	     �)  �X	     �)  �X	     *  �X	     +*  �X	     D*  �X	     X*  �X	     m*  �X	     �*  �X	     �*  �X	     �*  �X	     �*  �X	     �*  �X	     +  �X	     9+  �X	     ^+  �X	     +  �X	     �+  �X	     �+  �X	     �+  �X	     ,  �X	     2,   Y	     O,  Y	     q,  Y	     �,  Y	     �,  Y	     �,  Y	     �,  Y	     -  Y	     --   Y	     Q-  $Y	     t-  (Y	     �-  ,Y	     �-  0Y	     �-  4Y	     .  8Y	     ,.  <Y	     S.  @Y	     {.  DY	     �.  HY	     �.  LY	     �.  PY	     '/  TY	     G/  XY	     S2           ��`2  75U     y2  �[     �2  �[     �2  �[�    �2  �5Q     �2  �5S     3  06    3  17�     +3  �7�    Q3  C:e    {3  �<�    �3  K>R    �3  �?    �3  �@J     4  �@A    =4  -Ic    a4  �N�	    4  pXi     �4  �XC    �4  [�    �4  �g�    5  �p�    @5  ���    w5  s��    �5  4��    �5  ��    �#  �Y	     �#  �Y	     �#  �Y	     �#  �Y	     $  �Y	     2$  �Y	     C$  �Y	     T$  �Y	     e$  �Y	     |$  �Y	     �$  �Y	     �$  �Y	     �$  �Y	     �$  �Y	     �$  �Y	     %  �Y	     L%  �Y	     �%  �Y	     �%  �Y	     �%  �Y	     �%  �Y	     �%  �Y	     &   Z	     =&  Z	     i&  Z	     �&  Z	     �&  Z	     �&  Z	     �&  Z	     �&  Z	     )'   Z	     T'  $Z	     �'  (Z	     �'  ,Z	     �'  0Z	     (  4Z	     %(  8Z	     <(  <Z	     O(  @Z	     a(  DZ	     y(  HZ	     �(  LZ	     �(  PZ	     �(  TZ	     �(  XZ	     �(  \Z	     )  `Z	     )  dZ	     +)  hZ	     D)  lZ	     ])  pZ	     p)  tZ	     �)  xZ	     �)  |Z	     �)  �Z	     �)  �Z	     �)  �Z	     �)  �Z	     *  �Z	     +*  �Z	     D*  �Z	     X*  �Z	     m*  �Z	     �*  �Z	     �*  �Z	     �*  �Z	     �*  �Z	     �*  �Z	     +  �Z	     9+  �Z	     ^+  �Z	     +  �Z	     �+  �Z	     �+  �Z	     �+  �Z	     ,  �Z	     2,  �Z	     O,  �Z	     q,  �Z	     �,  �Z	     �,  �Z	     �,  �Z	     �,  �Z	     -  �Z	     --  �Z	     Q-  �Z	     t-   [	     �-  [	     �-  [	     �-  [	     .  [	     ,.  [	     S.  [	     {.  [	     �.   [	     �.  $[	     �.  ([	     '/  ,[	     G/  0[	     �5           ���#  8[	     �#  9[	     �#  :[	     �#  ;[	     $  <[	     2$  @[	     C$  D[	     T$  H[	     e$  L[	     |$  P[	     �$  T[	     �$  X[	     �$  \[	     �$  `[	     �$  d[	     %  h[	     L%  l[	     �%  p[	     �%  x[	     �%  |[	     �%  �[	     �%  �[	     &  �[	     =&  �[	     i&  �[	     �&  �[	     �&  �[	     �&  �[	     �&  �[	     �&  �[	     )'  �[	     T'  �[	     �'  �[	     �'  �[	     �'  �[	     (  �[	     %(  �[	     <(  �[	     O(  �[	     a(  �[	     y(  �[	     �(  �[	     �(  �[	     �(  �[	     �(  �[	     �(  �[	     )  �[	     )  �[	     +)  �[	     D)  �[	     ])  �[	     p)  �[	     �)   \	     �)  \	     �)  \	     �)  \	     �)  \	     �)  \	     *  \	     +*  \	     D*   \	     X*  $\	     m*  (\	     �*  ,\	     �*  0\	     �*  4\	     �*  8\	     �*  <\	     +  @\	     9+  D\	     ^+  H\	     +  L\	     �+  P\	     �+  T\	     �+  X\	     ,  \\	     2,  `\	     O,  d\	     q,  h\	     �,  l\	     �,  p\	     �,  t\	     �,  x\	     -  |\	     --  �\	     Q-  �\	     t-  �\	     �-  �\	     �-  �\	     �-  �\	     .  �\	     ,.  �\	     S.  �\	     {.  �\	     �.  �\	     �.  �\	     �.  �\	     '/  �\	     G/  �\	     �5           ���#  �\	     �#  �\	     �#  �\	     �#  �\	     $  �\	     2$  �\	     C$  �\	     T$  �\	     e$  �\	     |$  �\	     �$  �\	     �$  �\	     �$  �\	     �$  �\	     �$  �\	     %  �\	     L%  �\	     �%  �\	     �%   ]	     �%  ]	     �%  ]	     �%  ]	     &  ]	     =&  ]	     i&  ]	     �&  ]	     �&   ]	     �&  $]	     �&  (]	     �&  ,]	     )'  0]	     T'  4]	     �'  8]	     �'  <]	     �'  @]	     (  D]	     %(  H]	     <(  L]	     O(  P]	     a(  T]	     y(  X]	     �(  \]	     �(  `]	     �(  d]	     �(  h]	     �(  l]	     )  p]	     )  t]	     +)  x]	     D)  |]	     ])  �]	     p)  �]	     �)  �]	     �)  �]	     �)  �]	     �)  �]	     �)  �]	     �)  �]	     *  �]	     +*  �]	     D*  �]	     X*  �]	     m*  �]	     �*  �]	     �*  �]	     �*  �]	     �*  �]	     �*  �]	     +  �]	     9+  �]	     ^+  �]	     +  �]	     �+  �]	     �+  �]	     �+  �]	     ,  �]	     2,  �]	     O,  �]	     q,  �]	     �,  �]	     �,  �]	     �,  �]	     �,   ^	     -  ^	     --  ^	     Q-  ^	     t-  ^	     �-  ^	     �-  ^	     �-  ^	     .   ^	     ,.  $^	     S.  (^	     {.  ,^	     �.  0^	     �.  4^	     �.  8^	     '/  <^	     G/  @^	     6           ���#  H^	     �#  I^	     �#  J^	     �#  K^	     $  L^	     2$  P^	     C$  T^	     T$  X^	     e$  \^	     |$  `^	     �$  d^	     �$  h^	     �$  l^	     �$  p^	     �$  t^	     %  x^	     L%  |^	     �%  �^	     �%  �^	     �%  �^	     �%  �^	     �%  �^	     &  �^	     =&  �^	     i&  �^	     �&  �^	     �&  �^	     �&  �^	     �&  �^	     �&  �^	     )'  �^	     T'  �^	     �'  �^	     �'  �^	     �'  �^	     (  �^	     %(  �^	     <(  �^	     O(  �^	     a(  �^	     y(  �^	     �(  �^	     �(  �^	     �(  �^	     �(  �^	     �(  �^	     )  �^	     )  �^	     +)   _	     D)  _	     ])  _	     p)  _	     �)  _	     �)  _	     �)  _	     �)  _	     �)   _	     �)  $_	     *  (_	     +*  ,_	     D*  0_	     X*  4_	     m*  8_	     �*  <_	     �*  @_	     �*  D_	     �*  H_	     �*  L_	     +  P_	     9+  T_	     ^+  X_	     +  \_	     �+  `_	     �+  d_	     �+  h_	     ,  l_	     2,  p_	     O,  t_	     q,  x_	     �,  |_	     �,  �_	     �,  �_	     �,  �_	     -  �_	     --  �_	     Q-  �_	     t-  �_	     �-  �_	     �-  �_	     �-  �_	     .  �_	     ,.  �_	     S.  �_	     {.  �_	     �.  �_	     �.  �_	     �.  �_	     '/  �_	     G/  �_	     6           ���#  �_	     �#  �_	     �#  �_	     �#  �_	     $  �_	     2$  �_	     C$  �_	     T$  �_	     e$  �_	     |$  �_	     �$  �_	     �$  �_	     �$  �_	     �$  �_	     �$  �_	     %   `	     L%  `	     �%  `	     �%  `	     �%  `	     �%  `	     �%  `	     &   `	     =&  $`	     i&  (`	     �&  ,`	     �&  0`	     �&  4`	     �&  8`	     �&  <`	     )'  @`	     T'  D`	     �'  H`	     �'  L`	     �'  P`	     (  T`	     %(  X`	     <(  \`	     O(  ``	     a(  d`	     y(  h`	     �(  l`	     �(  p`	     �(  t`	     �(  x`	     �(  |`	     )  �`	     )  �`	     +)  �`	     D)  �`	     ])  �`	     p)  �`	     �)  �`	     �)  �`	     �)  �`	     �)  �`	     �)  �`	     �)  �`	     *  �`	     +*  �`	     D*  �`	     X*  �`	     m*  �`	     �*  �`	     �*  �`	     �*  �`	     �*  �`	     �*  �`	     +  �`	     9+  �`	     ^+  �`	     +  �`	     �+  �`	     �+  �`	     �+  �`	     ,  �`	     2,  �`	     O,  �`	     q,   a	     �,  a	     �,  a	     �,  a	     �,  a	     -  a	     --  a	     Q-  a	     t-   a	     �-  $a	     �-  (a	     �-  ,a	     .  0a	     ,.  4a	     S.  8a	     {.  <a	     �.  @a	     �.  Da	     �.  Ha	     '/  La	     G/  Pa	     %6           ���#  Xa	     �#  Ya	     �#  Za	     �#  [a	     $  \a	     2$  `a	     C$  da	     T$  ha	     e$  la	     |$  pa	     �$  ta	     �$  xa	     �$  |a	     �$  �a	     �$  �a	     %  �a	     L%  �a	     �%  �a	     �%  �a	     �%  �a	     �%  �a	     �%  �a	     &  �a	     =&  �a	     i&  �a	     �&  �a	     �&  �a	     �&  �a	     �&  �a	     �&  �a	     )'  �a	     T'  �a	     �'  �a	     �'  �a	     �'  �a	     (  �a	     %(  �a	     <(  �a	     O(  �a	     a(  �a	     y(  �a	     �(  �a	     �(  �a	     �(  �a	     �(   b	     �(  b	     )  b	     )  b	     +)  b	     D)  b	     ])  b	     p)  b	     �)   b	     �)  $b	     �)  (b	     �)  ,b	     �)  0b	     �)  4b	     *  8b	     +*  <b	     D*  @b	     X*  Db	     m*  Hb	     �*  Lb	     �*  Pb	     �*  Tb	     �*  Xb	     �*  \b	     +  `b	     9+  db	     ^+  hb	     +  lb	     �+  pb	     �+  tb	     �+  xb	     ,  |b	     2,  �b	     O,  �b	     q,  �b	     �,  �b	     �,  �b	     �,  �b	     �,  �b	     -  �b	     --  �b	     Q-  �b	     t-  �b	     �-  �b	     �-  �b	     �-  �b	     .  �b	     ,.  �b	     S.  �b	     {.  �b	     �.  �b	     �.  �b	     �.  �b	     '/  �b	     G/  �b	     B6           ���#  �b	     �#  �b	     �#  �b	     �#  �b	     $  �b	     2$  �b	     C$  �b	     T$  �b	     e$  �b	     |$  �b	     �$  �b	     �$   c	     �$  c	     �$  c	     �$  c	     %  c	     L%  c	     �%  c	     �%   c	     �%  $c	     �%  (c	     �%  ,c	     &  0c	     =&  4c	     i&  8c	     �&  <c	     �&  @c	     �&  Dc	     �&  Hc	     �&  Lc	     )'  Pc	     T'  Tc	     �'  Xc	     �'  \c	     �'  `c	     (  dc	     %(  hc	     <(  lc	     O(  pc	     a(  tc	     y(  xc	     �(  |c	     �(  �c	     �(  �c	     �(  �c	     �(  �c	     )  �c	     )  �c	     +)  �c	     D)  �c	     ])  �c	     p)  �c	     �)  �c	     �)  �c	     �)  �c	     �)  �c	     �)  �c	     �)  �c	     *  �c	     +*  �c	     D*  �c	     X*  �c	     m*  �c	     �*  �c	     �*  �c	     �*  �c	     �*  �c	     �*  �c	     +  �c	     9+  �c	     ^+  �c	     +  �c	     �+  �c	     �+  �c	     �+   d	     ,  d	     2,  d	     O,  d	     q,  d	     �,  d	     �,  d	     �,  d	     �,   d	     -  $d	     --  (d	     Q-  ,d	     t-  0d	     �-  4d	     �-  8d	     �-  <d	     .  @d	     ,.  Dd	     S.  Hd	     {.  Ld	     �.  Pd	     �.  Td	     �.  Xd	     '/  \d	     G/  `d	     M6           ���#  hd	     �#  id	     �#  jd	     �#  kd	     $  ld	     2$  pd	     C$  td	     T$  xd	     e$  |d	     |$  �d	     �$  �d	     �$  �d	     �$  �d	     �$  �d	     �$  �d	     %  �d	     L%  �d	     �%  �d	     �%  �d	     �%  �d	     �%  �d	     �%  �d	     &  �d	     =&  �d	     i&  �d	     �&  �d	     �&  �d	     �&  �d	     �&  �d	     �&  �d	     )'  �d	     T'  �d	     �'  �d	     �'  �d	     �'  �d	     (  �d	     %(  �d	     <(  �d	     O(  �d	     a(  �d	     y(   e	     �(  e	     �(  e	     �(  e	     �(  e	     �(  e	     )  e	     )  e	     +)   e	     D)  $e	     ])  (e	     p)  ,e	     �)  0e	     �)  4e	     �)  8e	     �)  <e	     �)  @e	     �)  De	     *  He	     +*  Le	     D*  Pe	     X*  Te	     m*  Xe	     �*  \e	     �*  `e	     �*  de	     �*  he	     �*  le	     +  pe	     9+  te	     ^+  xe	     +  |e	     �+  �e	     �+  �e	     �+  �e	     ,  �e	     2,  �e	     O,  �e	     q,  �e	     �,  �e	     �,  �e	     �,  �e	     �,  �e	     -  �e	     --  �e	     Q-  �e	     t-  �e	     �-  �e	     �-  �e	     �-  �e	     .  �e	     ,.  �e	     S.  �e	     {.  �e	     �.  �e	     �.  �e	     �.  �e	     '/  �e	     G/  �e	     a6           ���#  �e	     �#  �e	     �#  �e	     �#  �e	     $  �e	     2$  �e	     C$  �e	     T$   f	     e$  f	     |$  f	     �$  f	     �$  f	     �$  f	     �$  f	     �$  f	     %   f	     L%  $f	     �%  (f	     �%  0f	     �%  4f	     �%  8f	     �%  <f	     &  @f	     =&  Df	     i&  Hf	     �&  Lf	     �&  Pf	     �&  Tf	     �&  Xf	     �&  \f	     )'  `f	     T'  df	     �'  hf	     �'  lf	     �'  pf	     (  tf	     %(  xf	     <(  |f	     O(  �f	     a(  �f	     y(  �f	     �(  �f	     �(  �f	     �(  �f	     �(  �f	     �(  �f	     )  �f	     )  �f	     +)  �f	     D)  �f	     ])  �f	     p)  �f	     �)  �f	     �)  �f	     �)  �f	     �)  �f	     �)  �f	     �)  �f	     *  �f	     +*  �f	     D*  �f	     X*  �f	     m*  �f	     �*  �f	     �*  �f	     �*  �f	     �*  �f	     �*  �f	     +  �f	     9+  �f	     ^+   g	     +  g	     �+  g	     �+  g	     �+  g	     ,  g	     2,  g	     O,  g	     q,   g	     �,  $g	     �,  (g	     �,  ,g	     �,  0g	     -  4g	     --  8g	     Q-  <g	     t-  @g	     �-  Dg	     �-  Hg	     �-  Lg	     .  Pg	     ,.  Tg	     S.  Xg	     {.  \g	     �.  `g	     �.  dg	     �.  hg	     '/  lg	     G/  pg	     l6           ���#  xg	     �#  yg	     �#  zg	     �#  {g	     $  |g	     2$  �g	     C$  �g	     T$  �g	     e$  �g	     |$  �g	     �$  �g	     �$  �g	     �$  �g	     �$  �g	     �$  �g	     %  �g	     L%  �g	     �%  �g	     �%  �g	     �%  �g	     �%  �g	     �%  �g	     &  �g	     =&  �g	     i&  �g	     �&  �g	     �&  �g	     �&  �g	     �&  �g	     �&  �g	     )'  �g	     T'  �g	     �'  �g	     �'  �g	     �'  �g	     (  �g	     %(   h	     <(  h	     O(  h	     a(  h	     y(  h	     �(  h	     �(  h	     �(  h	     �(   h	     �(  $h	     )  (h	     )  ,h	     +)  0h	     D)  4h	     ])  8h	     p)  <h	     �)  @h	     �)  Dh	     �)  Hh	     �)  Lh	     �)  Ph	     �)  Th	     *  Xh	     +*  \h	     D*  `h	     X*  dh	     m*  hh	     �*  lh	     �*  ph	     �*  th	     �*  xh	     �*  |h	     +  �h	     9+  �h	     ^+  �h	     +  �h	     �+  �h	     �+  �h	     �+  �h	     ,  �h	     2,  �h	     O,  �h	     q,  �h	     �,  �h	     �,  �h	     �,  �h	     �,  �h	     -  �h	     --  �h	     Q-  �h	     t-  �h	     �-  �h	     �-  �h	     �-  �h	     .  �h	     ,.  �h	     S.  �h	     {.  �h	     �.  �h	     �.  �h	     �.  �h	     '/  �h	     G/  �h	     �6           ���#   i	     �#  i	     �#  i	     �#  i	     $  i	     2$  i	     C$  i	     T$  i	     e$  i	     |$  i	     �$  i	     �$   i	     �$  $i	     �$  (i	     �$  ,i	     %  0i	     L%  4i	     �%  8i	     �%  @i	     �%  Di	     �%  Hi	     �%  Li	     &  Pi	     =&  Ti	     i&  Xi	     �&  \i	     �&  `i	     �&  di	     �&  hi	     �&  li	     )'  pi	     T'  ti	     �'  xi	     �'  |i	     �'  �i	     (  �i	     %(  �i	     <(  �i	     O(  �i	     a(  �i	     y(  �i	     �(  �i	     �(  �i	     �(  �i	     �(  �i	     �(  �i	     )  �i	     )  �i	     +)  �i	     D)  �i	     ])  �i	     p)  �i	     �)  �i	     �)  �i	     �)  �i	     �)  �i	     �)  �i	     �)  �i	     *  �i	     +*  �i	     D*  �i	     X*  �i	     m*  �i	     �*  �i	     �*  �i	     �*  �i	     �*   j	     �*  j	     +  j	     9+  j	     ^+  j	     +  j	     �+  j	     �+  j	     �+   j	     ,  $j	     2,  (j	     O,  ,j	     q,  0j	     �,  4j	     �,  8j	     �,  <j	     �,  @j	     -  Dj	     --  Hj	     Q-  Lj	     t-  Pj	     �-  Tj	     �-  Xj	     �-  \j	     .  `j	     ,.  dj	     S.  hj	     {.  lj	     �.  pj	     �.  tj	     �.  xj	     '/  |j	     G/  �j	     �6           ���#  �j	     �#  �j	     �#  �j	     �#  �j	     $  �j	     2$  �j	     C$  �j	     T$  �j	     e$  �j	     |$  �j	     �$  �j	     �$  �j	     �$  �j	     �$  �j	     �$  �j	     %  �j	     L%  �j	     �%  �j	     �%  �j	     �%  �j	     �%  �j	     �%  �j	     &  �j	     =&  �j	     i&  �j	     �&  �j	     �&  �j	     �&  �j	     �&  �j	     �&  �j	     )'  �j	     T'  �j	     �'   k	     �'  k	     �'  k	     (  k	     %(  k	     <(  k	     O(  k	     a(  k	     y(   k	     �(  $k	     �(  (k	     �(  ,k	     �(  0k	     �(  4k	     )  8k	     )  <k	     +)  @k	     D)  Dk	     ])  Hk	     p)  Lk	     �)  Pk	     �)  Tk	     �)  Xk	     �)  \k	     �)  `k	     �)  dk	     *  hk	     +*  lk	     D*  pk	     X*  tk	     m*  xk	     �*  |k	     �*  �k	     �*  �k	     �*  �k	     �*  �k	     +  �k	     9+  �k	     ^+  �k	     +  �k	     �+  �k	     �+  �k	     �+  �k	     ,  �k	     2,  �k	     O,  �k	     q,  �k	     �,  �k	     �,  �k	     �,  �k	     �,  �k	     -  �k	     --  �k	     Q-  �k	     t-  �k	     �-  �k	     �-  �k	     �-  �k	     .  �k	     ,.  �k	     S.  �k	     {.  �k	     �.  �k	     �.  �k	     �.   l	     '/  l	     G/  l	     �6           ���#  l	     �#  l	     �#  l	     �#  l	     $  l	     2$  l	     C$  l	     T$   l	     e$  $l	     |$  (l	     �$  ,l	     �$  0l	     �$  4l	     �$  8l	     �$  <l	     %  @l	     L%  Dl	     �%  Hl	     �%  Pl	     �%  Tl	     �%  Xl	     �%  \l	     &  `l	     =&  dl	     i&  hl	     �&  ll	     �&  pl	     �&  tl	     �&  xl	     �&  |l	     )'  �l	     T'  �l	     �'  �l	     �'  �l	     �'  �l	     (  �l	     %(  �l	     <(  �l	     O(  �l	     a(  �l	     y(  �l	     �(  �l	     �(  �l	     �(  �l	     �(  �l	     �(  �l	     )  �l	     )  �l	     +)  �l	     D)  �l	     ])  �l	     p)  �l	     �)  �l	     �)  �l	     �)  �l	     �)  �l	     �)  �l	     �)  �l	     *  �l	     +*  �l	     D*  �l	     X*  �l	     m*   m	     �*  m	     �*  m	     �*  m	     �*  m	     �*  m	     +  m	     9+  m	     ^+   m	     +  $m	     �+  (m	     �+  ,m	     �+  0m	     ,  4m	     2,  8m	     O,  <m	     q,  @m	     �,  Dm	     �,  Hm	     �,  Lm	     �,  Pm	     -  Tm	     --  Xm	     Q-  \m	     t-  `m	     �-  dm	     �-  hm	     �-  lm	     .  pm	     ,.  tm	     S.  xm	     {.  |m	     �.  �m	     �.  �m	     �.  �m	     '/  �m	     G/  �m	     �6           ���#  �m	     �#  �m	     �#  �m	     �#  �m	     $  �m	     2$  �m	     C$  �m	     T$  �m	     e$  �m	     |$  �m	     �$  �m	     �$  �m	     �$  �m	     �$  �m	     �$  �m	     %  �m	     L%  �m	     �%  �m	     �%  �m	     �%  �m	     �%  �m	     �%  �m	     &  �m	     =&  �m	     i&  �m	     �&  �m	     �&  �m	     �&  �m	     �&   n	     �&  n	     )'  n	     T'  n	     �'  n	     �'  n	     �'  n	     (  n	     %(   n	     <(  $n	     O(  (n	     a(  ,n	     y(  0n	     �(  4n	     �(  8n	     �(  <n	     �(  @n	     �(  Dn	     )  Hn	     )  Ln	     +)  Pn	     D)  Tn	     ])  Xn	     p)  \n	     �)  `n	     �)  dn	     �)  hn	     �)  ln	     �)  pn	     �)  tn	     *  xn	     +*  |n	     D*  �n	     X*  �n	     m*  �n	     �*  �n	     �*  �n	     �*  �n	     �*  �n	     �*  �n	     +  �n	     9+  �n	     ^+  �n	     +  �n	     �+  �n	     �+  �n	     �+  �n	     ,  �n	     2,  �n	     O,  �n	     q,  �n	     �,  �n	     �,  �n	     �,  �n	     �,  �n	     -  �n	     --  �n	     Q-  �n	     t-  �n	     �-  �n	     �-  �n	     �-  �n	     .  �n	     ,.  �n	     S.   o	     {.  o	     �.  o	     �.  o	     �.  o	     '/  o	     G/  o	     �6           ���#   o	     �#  !o	     �#  "o	     �#  #o	     $  $o	     2$  (o	     C$  ,o	     T$  0o	     e$  4o	     |$  8o	     �$  <o	     �$  @o	     �$  Do	     �$  Ho	     �$  Lo	     %  Po	     L%  To	     �%  Xo	     �%  `o	     �%  do	     �%  ho	     �%  lo	     &  po	     =&  to	     i&  xo	     �&  |o	     �&  �o	     �&  �o	     �&  �o	     �&  �o	     )'  �o	     T'  �o	     �'  �o	     �'  �o	     �'  �o	     (  �o	     %(  �o	     <(  �o	     O(  �o	     a(  �o	     y(  �o	     �(  �o	     �(  �o	     �(  �o	     �(  �o	     �(  �o	     )  �o	     )  �o	     +)  �o	     D)  �o	     ])  �o	     p)  �o	     �)  �o	     �)  �o	     �)  �o	     �)  �o	     �)  �o	     �)  �o	     *   p	     +*  p	     D*  p	     X*  p	     m*  p	     �*  p	     �*  p	     �*  p	     �*   p	     �*  $p	     +  (p	     9+  ,p	     ^+  0p	     +  4p	     �+  8p	     �+  <p	     �+  @p	     ,  Dp	     2,  Hp	     O,  Lp	     q,  Pp	     �,  Tp	     �,  Xp	     �,  \p	     �,  `p	     -  dp	     --  hp	     Q-  lp	     t-  pp	     �-  tp	     �-  xp	     �-  |p	     .  �p	     ,.  �p	     S.  �p	     {.  �p	     �.  �p	     �.  �p	     �.  �p	     '/  �p	     G/  �p	     �6           ���#  �p	     �#  �p	     �#  �p	     �#  �p	     $  �p	     2$  �p	     C$  �p	     T$  �p	     e$  �p	     |$  �p	     �$  �p	     �$  �p	     �$  �p	     �$  �p	     �$  �p	     %  �p	     L%  �p	     �%  �p	     �%  �p	     �%  �p	     �%  �p	     �%  �p	     &  �p	     =&  �p	     i&   q	     �&  q	     �&  q	     �&  q	     �&  q	     �&  q	     )'  q	     T'  q	     �'   q	     �'  $q	     �'  (q	     (  ,q	     %(  0q	     <(  4q	     O(  8q	     a(  <q	     y(  @q	     �(  Dq	     �(  Hq	     �(  Lq	     �(  Pq	     �(  Tq	     )  Xq	     )  \q	     +)  `q	     D)  dq	     ])  hq	     p)  lq	     �)  pq	     �)  tq	     �)  xq	     �)  |q	     �)  �q	     �)  �q	     *  �q	     +*  �q	     D*  �q	     X*  �q	     m*  �q	     �*  �q	     �*  �q	     �*  �q	     �*  �q	     �*  �q	     +  �q	     9+  �q	     ^+  �q	     +  �q	     �+  �q	     �+  �q	     �+  �q	     ,  �q	     2,  �q	     O,  �q	     q,  �q	     �,  �q	     �,  �q	     �,  �q	     �,  �q	     -  �q	     --  �q	     Q-  �q	     t-  �q	     �-  �q	     �-   r	     �-  r	     .  r	     ,.  r	     S.  r	     {.  r	     �.  r	     �.  r	     �.   r	     '/  $r	     G/  (r	     �6           ���#  0r	     �#  1r	     �#  2r	     �#  3r	     $  4r	     2$  8r	     C$  <r	     T$  @r	     e$  Dr	     |$  Hr	     �$  Lr	     �$  Pr	     �$  Tr	     �$  Xr	     �$  \r	     %  `r	     L%  dr	     �%  hr	     �%  pr	     �%  tr	     �%  xr	     �%  |r	     &  �r	     =&  �r	     i&  �r	     �&  �r	     �&  �r	     �&  �r	     �&  �r	     �&  �r	     )'  �r	     T'  �r	     �'  �r	     �'  �r	     �'  �r	     (  �r	     %(  �r	     <(  �r	     O(  �r	     a(  �r	     y(  �r	     �(  �r	     �(  �r	     �(  �r	     �(  �r	     �(  �r	     )  �r	     )  �r	     +)  �r	     D)  �r	     ])  �r	     p)  �r	     �)  �r	     �)  �r	     �)   s	     �)  s	     �)  s	     �)  s	     *  s	     +*  s	     D*  s	     X*  s	     m*   s	     �*  $s	     �*  (s	     �*  ,s	     �*  0s	     �*  4s	     +  8s	     9+  <s	     ^+  @s	     +  Ds	     �+  Hs	     �+  Ls	     �+  Ps	     ,  Ts	     2,  Xs	     O,  \s	     q,  `s	     �,  ds	     �,  hs	     �,  ls	     �,  ps	     -  ts	     --  xs	     Q-  |s	     t-  �s	     �-  �s	     �-  �s	     �-  �s	     .  �s	     ,.  �s	     S.  �s	     {.  �s	     �.  �s	     �.  �s	     �.  �s	     '/  �s	     G/  �s	     �6           ���#  �s	     �#  �s	     �#  �s	     �#  �s	     $  �s	     2$  �s	     C$  �s	     T$  �s	     e$  �s	     |$  �s	     �$  �s	     �$  �s	     �$  �s	     �$  �s	     �$  �s	     %  �s	     L%  �s	     �%  �s	     �%  �s	     �%  �s	     �%   t	     �%  t	     &  t	     =&  t	     i&  t	     �&  t	     �&  t	     �&  t	     �&   t	     �&  $t	     )'  (t	     T'  ,t	     �'  0t	     �'  4t	     �'  8t	     (  <t	     %(  @t	     <(  Dt	     O(  Ht	     a(  Lt	     y(  Pt	     �(  Tt	     �(  Xt	     �(  \t	     �(  `t	     �(  dt	     )  ht	     )  lt	     +)  pt	     D)  tt	     ])  xt	     p)  |t	     �)  �t	     �)  �t	     �)  �t	     �)  �t	     �)  �t	     �)  �t	     *  �t	     +*  �t	     D*  �t	     X*  �t	     m*  �t	     �*  �t	     �*  �t	     �*  �t	     �*  �t	     �*  �t	     +  �t	     9+  �t	     ^+  �t	     +  �t	     �+  �t	     �+  �t	     �+  �t	     ,  �t	     2,  �t	     O,  �t	     q,  �t	     �,  �t	     �,  �t	     �,  �t	     �,  �t	     -  �t	     --   u	     Q-  u	     t-  u	     �-  u	     �-  u	     �-  u	     .  u	     ,.  u	     S.   u	     {.  $u	     �.  (u	     �.  ,u	     �.  0u	     '/  4u	     G/  8u	     �6           ���#  @u	     �#  Au	     �#  Bu	     �#  Cu	     $  Du	     2$  Hu	     C$  Lu	     T$  Pu	     e$  Tu	     |$  Xu	     �$  \u	     �$  `u	     �$  du	     �$  hu	     �$  lu	     %  pu	     L%  tu	     �%  xu	     �%  �u	     �%  �u	     �%  �u	     �%  �u	     &  �u	     =&  �u	     i&  �u	     �&  �u	     �&  �u	     �&  �u	     �&  �u	     �&  �u	     )'  �u	     T'  �u	     �'  �u	     �'  �u	     �'  �u	     (  �u	     %(  �u	     <(  �u	     O(  �u	     a(  �u	     y(  �u	     �(  �u	     �(  �u	     �(  �u	     �(  �u	     �(  �u	     )  �u	     )  �u	     +)  �u	     D)  �u	     ])   v	     p)  v	     �)  v	     �)  v	     �)  v	     �)  v	     �)  v	     �)  v	     *   v	     +*  $v	     D*  (v	     X*  ,v	     m*  0v	     �*  4v	     �*  8v	     �*  <v	     �*  @v	     �*  Dv	     +  Hv	     9+  Lv	     ^+  Pv	     +  Tv	     �+  Xv	     �+  \v	     �+  `v	     ,  dv	     2,  hv	     O,  lv	     q,  pv	     �,  tv	     �,  xv	     �,  |v	     �,  �v	     -  �v	     --  �v	     Q-  �v	     t-  �v	     �-  �v	     �-  �v	     �-  �v	     .  �v	     ,.  �v	     S.  �v	     {.  �v	     �.  �v	     �.  �v	     �.  �v	     '/  �v	     G/  �v	     7           ���#  �v	     �#  �v	     �#  �v	     �#  �v	     $  �v	     2$  �v	     C$  �v	     T$  �v	     e$  �v	     |$  �v	     �$  �v	     �$  �v	     �$  �v	     �$  �v	     �$  �v	     %  �v	     L%  �v	     �%   w	     �%  w	     �%  w	     �%  w	     �%  w	     &  w	     =&  w	     i&   w	     �&  $w	     �&  (w	     �&  ,w	     �&  0w	     �&  4w	     )'  8w	     T'  <w	     �'  @w	     �'  Dw	     �'  Hw	     (  Lw	     %(  Pw	     <(  Tw	     O(  Xw	     a(  \w	     y(  `w	     �(  dw	     �(  hw	     �(  lw	     �(  pw	     �(  tw	     )  xw	     )  |w	     +)  �w	     D)  �w	     ])  �w	     p)  �w	     �)  �w	     �)  �w	     �)  �w	     �)  �w	     �)  �w	     �)  �w	     *  �w	     +*  �w	     D*  �w	     X*  �w	     m*  �w	     �*  �w	     �*  �w	     �*  �w	     �*  �w	     �*  �w	     +  �w	     9+  �w	     ^+  �w	     +  �w	     �+  �w	     �+  �w	     �+  �w	     ,  �w	     2,  �w	     O,  �w	     q,  �w	     �,  �w	     �,   x	     �,  x	     �,  x	     -  x	     --  x	     Q-  x	     t-  x	     �-  x	     �-   x	     �-  $x	     .  (x	     ,.  ,x	     S.  0x	     {.  4x	     �.  8x	     �.  <x	     �.  @x	     '/  Dx	     G/  Hx	     7           ���#  Px	     �#  Qx	     �#  Rx	     �#  Sx	     $  Tx	     2$  Xx	     C$  \x	     T$  `x	     e$  dx	     |$  hx	     �$  lx	     �$  px	     �$  tx	     �$  xx	     �$  |x	     %  �x	     L%  �x	     �%  �x	     �%  �x	     �%  �x	     �%  �x	     �%  �x	     &  �x	     =&  �x	     i&  �x	     �&  �x	     �&  �x	     �&  �x	     �&  �x	     �&  �x	     )'  �x	     T'  �x	     �'  �x	     �'  �x	     �'  �x	     (  �x	     %(  �x	     <(  �x	     O(  �x	     a(  �x	     y(  �x	     �(  �x	     �(  �x	     �(  �x	     �(  �x	     �(  �x	     )   y	     )  y	     +)  y	     D)  y	     ])  y	     p)  y	     �)  y	     �)  y	     �)   y	     �)  $y	     �)  (y	     �)  ,y	     *  0y	     +*  4y	     D*  8y	     X*  <y	     m*  @y	     �*  Dy	     �*  Hy	     �*  Ly	     �*  Py	     �*  Ty	     +  Xy	     9+  \y	     ^+  `y	     +  dy	     �+  hy	     �+  ly	     �+  py	     ,  ty	     2,  xy	     O,  |y	     q,  �y	     �,  �y	     �,  �y	     �,  �y	     �,  �y	     -  �y	     --  �y	     Q-  �y	     t-  �y	     �-  �y	     �-  �y	     �-  �y	     .  �y	     ,.  �y	     S.  �y	     {.  �y	     �.  �y	     �.  �y	     �.  �y	     '/  �y	     G/  �y	     $7           ���#  �y	     �#  �y	     �#  �y	     �#  �y	     $  �y	     2$  �y	     C$  �y	     T$  �y	     e$  �y	     |$  �y	     �$  �y	     �$  �y	     �$  �y	     �$   z	     �$  z	     %  z	     L%  z	     �%  z	     �%  z	     �%  z	     �%   z	     �%  $z	     &  (z	     =&  ,z	     i&  0z	     �&  4z	     �&  8z	     �&  <z	     �&  @z	     �&  Dz	     )'  Hz	     T'  Lz	     �'  Pz	     �'  Tz	     �'  Xz	     (  \z	     %(  `z	     <(  dz	     O(  hz	     a(  lz	     y(  pz	     �(  tz	     �(  xz	     �(  |z	     �(  �z	     �(  �z	     )  �z	     )  �z	     +)  �z	     D)  �z	     ])  �z	     p)  �z	     �)  �z	     �)  �z	     �)  �z	     �)  �z	     �)  �z	     �)  �z	     *  �z	     +*  �z	     D*  �z	     X*  �z	     m*  �z	     �*  �z	     �*  �z	     �*  �z	     �*  �z	     �*  �z	     +  �z	     9+  �z	     ^+  �z	     +  �z	     �+  �z	     �+  �z	     �+  �z	     ,  �z	     2,   {	     O,  {	     q,  {	     �,  {	     �,  {	     �,  {	     �,  {	     -  {	     --   {	     Q-  ${	     t-  ({	     �-  ,{	     �-  0{	     �-  4{	     .  8{	     ,.  <{	     S.  @{	     {.  D{	     �.  H{	     �.  L{	     �.  P{	     '/  T{	     G/  X{	     :7           ���#  `{	     �#  a{	     �#  b{	     �#  c{	     $  d{	     2$  h{	     C$  l{	     T$  p{	     e$  t{	     |$  x{	     �$  |{	     �$  �{	     �$  �{	     �$  �{	     �$  �{	     %  �{	     L%  �{	     �%  �{	     �%  �{	     �%  �{	     �%  �{	     �%  �{	     &  �{	     =&  �{	     i&  �{	     �&  �{	     �&  �{	     �&  �{	     �&  �{	     �&  �{	     )'  �{	     T'  �{	     �'  �{	     �'  �{	     �'  �{	     (  �{	     %(  �{	     <(  �{	     O(  �{	     a(  �{	     y(  �{	     �(  �{	     �(   |	     �(  |	     �(  |	     �(  |	     )  |	     )  |	     +)  |	     D)  |	     ])   |	     p)  $|	     �)  (|	     �)  ,|	     �)  0|	     �)  4|	     �)  8|	     �)  <|	     *  @|	     +*  D|	     D*  H|	     X*  L|	     m*  P|	     �*  T|	     �*  X|	     �*  \|	     �*  `|	     �*  d|	     +  h|	     9+  l|	     ^+  p|	     +  t|	     �+  x|	     �+  ||	     �+  �|	     ,  �|	     2,  �|	     O,  �|	     q,  �|	     �,  �|	     �,  �|	     �,  �|	     �,  �|	     -  �|	     --  �|	     Q-  �|	     t-  �|	     �-  �|	     �-  �|	     �-  �|	     .  �|	     ,.  �|	     S.  �|	     {.  �|	     �.  �|	     �.  �|	     �.  �|	     '/  �|	     G/  �|	     D7           ���#  �|	     �#  �|	     �#  �|	     �#  �|	     $  �|	     2$  �|	     C$  �|	     T$  �|	     e$  �|	     |$   }	     �$  }	     �$  }	     �$  }	     �$  }	     �$  }	     %  }	     L%  }	     �%   }	     �%  (}	     �%  ,}	     �%  0}	     �%  4}	     &  8}	     =&  <}	     i&  @}	     �&  D}	     �&  H}	     �&  L}	     �&  P}	     �&  T}	     )'  X}	     T'  \}	     �'  `}	     �'  d}	     �'  h}	     (  l}	     %(  p}	     <(  t}	     O(  x}	     a(  |}	     y(  �}	     �(  �}	     �(  �}	     �(  �}	     �(  �}	     �(  �}	     )  �}	     )  �}	     +)  �}	     D)  �}	     ])  �}	     p)  �}	     �)  �}	     �)  �}	     �)  �}	     �)  �}	     �)  �}	     �)  �}	     *  �}	     +*  �}	     D*  �}	     X*  �}	     m*  �}	     �*  �}	     �*  �}	     �*  �}	     �*  �}	     �*  �}	     +  �}	     9+  �}	     ^+  �}	     +  �}	     �+   ~	     �+  ~	     �+  ~	     ,  ~	     2,  ~	     O,  ~	     q,  ~	     �,  ~	     �,   ~	     �,  $~	     �,  (~	     -  ,~	     --  0~	     Q-  4~	     t-  8~	     �-  <~	     �-  @~	     �-  D~	     .  H~	     ,.  L~	     S.  P~	     {.  T~	     �.  X~	     �.  \~	     �.  `~	     '/  d~	     G/  h~	     Z7           ���#  p~	     �#  q~	     �#  r~	     �#  s~	     $  t~	     2$  x~	     C$  |~	     T$  �~	     e$  �~	     |$  �~	     �$  �~	     �$  �~	     �$  �~	     �$  �~	     �$  �~	     %  �~	     L%  �~	     �%  �~	     �%  �~	     �%  �~	     �%  �~	     �%  �~	     &  �~	     =&  �~	     i&  �~	     �&  �~	     �&  �~	     �&  �~	     �&  �~	     �&  �~	     )'  �~	     T'  �~	     �'  �~	     �'  �~	     �'  �~	     (  �~	     %(  �~	     <(  �~	     O(   	     a(  	     y(  	     �(  	     �(  	     �(  	     �(  	     �(  	     )   	     )  $	     +)  (	     D)  ,	     ])  0	     p)  4	     �)  8	     �)  <	     �)  @	     �)  D	     �)  H	     �)  L	     *  P	     +*  T	     D*  X	     X*  \	     m*  `	     �*  d	     �*  h	     �*  l	     �*  p	     �*  t	     +  x	     9+  |	     ^+  �	     +  �	     �+  �	     �+  �	     �+  �	     ,  �	     2,  �	     O,  �	     q,  �	     �,  �	     �,  �	     �,  �	     �,  �	     -  �	     --  �	     Q-  �	     t-  �	     �-  �	     �-  �	     �-  �	     .  �	     ,.  �	     S.  �	     {.  �	     �.  �	     �.  �	     �.  �	     '/  �	     G/  �	     e7           ���#  �	     �#  �	     �#  �	     �#  �	     $  �	     2$   �	     C$  �	     T$  �	     e$  �	     |$  �	     �$  �	     �$  �	     �$  �	     �$   �	     �$  $�	     %  (�	     L%  ,�	     �%  0�	     �%  8�	     �%  <�	     �%  @�	     �%  D�	     &  H�	     =&  L�	     i&  P�	     �&  T�	     �&  X�	     �&  \�	     �&  `�	     �&  d�	     )'  h�	     T'  l�	     �'  p�	     �'  t�	     �'  x�	     (  |�	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  Ā	     �)  Ȁ	     �)  ̀	     �)  Ѐ	     �)  Ԁ	     *  ؀	     +*  ܀	     D*  ��	     X*  �	     m*  �	     �*  �	     �*  ��	     �*  �	     �*  ��	     �*  ��	     +   �	     9+  �	     ^+  �	     +  �	     �+  �	     �+  �	     �+  �	     ,  �	     2,   �	     O,  $�	     q,  (�	     �,  ,�	     �,  0�	     �,  4�	     �,  8�	     -  <�	     --  @�	     Q-  D�	     t-  H�	     �-  L�	     �-  P�	     �-  T�	     .  X�	     ,.  \�	     S.  `�	     {.  d�	     �.  h�	     �.  l�	     �.  p�	     '/  t�	     G/  x�	     {7           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ā	     �%  ȁ	     �%  ́	     &  Ё	     =&  ԁ	     i&  ؁	     �&  ܁	     �&  ��	     �&  �	     �&  �	     �&  �	     )'  ��	     T'  �	     �'  ��	     �'  ��	     �'   �	     (  �	     %(  �	     <(  �	     O(  �	     a(  �	     y(  �	     �(  �	     �(   �	     �(  $�	     �(  (�	     �(  ,�	     )  0�	     )  4�	     +)  8�	     D)  <�	     ])  @�	     p)  D�	     �)  H�	     �)  L�	     �)  P�	     �)  T�	     �)  X�	     �)  \�	     *  `�	     +*  d�	     D*  h�	     X*  l�	     m*  p�	     �*  t�	     �*  x�	     �*  |�	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  Ă	     --  Ȃ	     Q-  ̂	     t-  Ђ	     �-  Ԃ	     �-  ؂	     �-  ܂	     .  ��	     ,.  �	     S.  �	     {.  �	     �.  ��	     �.  �	     �.  ��	     '/  ��	     G/   �	     �7           ���#  �	     �#  	�	     �#  
�	     �#  �	     $  �	     2$  �	     C$  �	     T$  �	     e$  �	     |$   �	     �$  $�	     �$  (�	     �$  ,�	     �$  0�	     �$  4�	     %  8�	     L%  <�	     �%  @�	     �%  H�	     �%  L�	     �%  P�	     �%  T�	     &  X�	     =&  \�	     i&  `�	     �&  d�	     �&  h�	     �&  l�	     �&  p�	     �&  t�	     )'  x�	     T'  |�	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ă	     ])  ȃ	     p)  ̃	     �)  Ѓ	     �)  ԃ	     �)  ؃	     �)  ܃	     �)  ��	     �)  �	     *  �	     +*  �	     D*  ��	     X*  �	     m*  ��	     �*  ��	     �*   �	     �*  �	     �*  �	     �*  �	     +  �	     9+  �	     ^+  �	     +  �	     �+   �	     �+  $�	     �+  (�	     ,  ,�	     2,  0�	     O,  4�	     q,  8�	     �,  <�	     �,  @�	     �,  D�	     �,  H�	     -  L�	     --  P�	     Q-  T�	     t-  X�	     �-  \�	     �-  `�	     �-  d�	     .  h�	     ,.  l�	     S.  p�	     {.  t�	     �.  x�	     �.  |�	     �.  ��	     '/  ��	     G/  ��	     �7           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  Ą	     �%  Ȅ	     �%  Є	     �%  Ԅ	     �%  ؄	     �%  ܄	     &  ��	     =&  �	     i&  �	     �&  �	     �&  ��	     �&  �	     �&  ��	     �&  ��	     )'   �	     T'  �	     �'  �	     �'  �	     �'  �	     (  �	     %(  �	     <(  �	     O(   �	     a(  $�	     y(  (�	     �(  ,�	     �(  0�	     �(  4�	     �(  8�	     �(  <�	     )  @�	     )  D�	     +)  H�	     D)  L�	     ])  P�	     p)  T�	     �)  X�	     �)  \�	     �)  `�	     �)  d�	     �)  h�	     �)  l�	     *  p�	     +*  t�	     D*  x�	     X*  |�	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ą	     �,  ȅ	     �,  ̅	     �,  Ѕ	     -  ԅ	     --  ؅	     Q-  ܅	     t-  ��	     �-  �	     �-  �	     �-  �	     .  ��	     ,.  �	     S.  ��	     {.  ��	     �.   �	     �.  �	     �.  �	     '/  �	     G/  �	     �7           ���#  �	     �#  �	     �#  �	     �#  �	     $  �	     2$   �	     C$  $�	     T$  (�	     e$  ,�	     |$  0�	     �$  4�	     �$  8�	     �$  <�	     �$  @�	     �$  D�	     %  H�	     L%  L�	     �%  P�	     �%  X�	     �%  \�	     �%  `�	     �%  d�	     &  h�	     =&  l�	     i&  p�	     �&  t�	     �&  x�	     �&  |�	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  Ć	     )  Ȇ	     )  ̆	     +)  І	     D)  Ԇ	     ])  ؆	     p)  ܆	     �)  ��	     �)  �	     �)  �	     �)  �	     �)  ��	     �)  �	     *  ��	     +*  ��	     D*   �	     X*  �	     m*  �	     �*  �	     �*  �	     �*  �	     �*  �	     �*  �	     +   �	     9+  $�	     ^+  (�	     +  ,�	     �+  0�	     �+  4�	     �+  8�	     ,  <�	     2,  @�	     O,  D�	     q,  H�	     �,  L�	     �,  P�	     �,  T�	     �,  X�	     -  \�	     --  `�	     Q-  d�	     t-  h�	     �-  l�	     �-  p�	     �-  t�	     .  x�	     ,.  |�	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �7           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ć	     �$  ȇ	     �$  ̇	     %  Ї	     L%  ԇ	     �%  ؇	     �%  ��	     �%  �	     �%  �	     �%  �	     &  ��	     =&  �	     i&  ��	     �&  ��	     �&   �	     �&  �	     �&  �	     �&  �	     )'  �	     T'  �	     �'  �	     �'  �	     �'   �	     (  $�	     %(  (�	     <(  ,�	     O(  0�	     a(  4�	     y(  8�	     �(  <�	     �(  @�	     �(  D�	     �(  H�	     �(  L�	     )  P�	     )  T�	     +)  X�	     D)  \�	     ])  `�	     p)  d�	     �)  h�	     �)  l�	     �)  p�	     �)  t�	     �)  x�	     �)  |�	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  Ĉ	     2,  Ȉ	     O,  ̈	     q,  Ј	     �,  Ԉ	     �,  ؈	     �,  ܈	     �,  ��	     -  �	     --  �	     Q-  �	     t-  ��	     �-  �	     �-  ��	     �-  ��	     .   �	     ,.  �	     S.  �	     {.  �	     �.  �	     �.  �	     �.  �	     '/  �	     G/   �	     �7           ���#  (�	     �#  )�	     �#  *�	     �#  +�	     $  ,�	     2$  0�	     C$  4�	     T$  8�	     e$  <�	     |$  @�	     �$  D�	     �$  H�	     �$  L�	     �$  P�	     �$  T�	     %  X�	     L%  \�	     �%  `�	     �%  h�	     �%  l�	     �%  p�	     �%  t�	     &  x�	     =&  |�	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ĉ	     �(  ȉ	     �(  ̉	     �(  Љ	     �(  ԉ	     )  ؉	     )  ܉	     +)  ��	     D)  �	     ])  �	     p)  �	     �)  ��	     �)  �	     �)  ��	     �)  ��	     �)   �	     �)  �	     *  �	     +*  �	     D*  �	     X*  �	     m*  �	     �*  �	     �*   �	     �*  $�	     �*  (�	     �*  ,�	     +  0�	     9+  4�	     ^+  8�	     +  <�	     �+  @�	     �+  D�	     �+  H�	     ,  L�	     2,  P�	     O,  T�	     q,  X�	     �,  \�	     �,  `�	     �,  d�	     �,  h�	     -  l�	     --  p�	     Q-  t�	     t-  x�	     �-  |�	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �7           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  Ċ	     |$  Ȋ	     �$  ̊	     �$  Њ	     �$  Ԋ	     �$  ؊	     �$  ܊	     %  ��	     L%  �	     �%  �	     �%  ��	     �%  �	     �%  ��	     �%  ��	     &   �	     =&  �	     i&  �	     �&  �	     �&  �	     �&  �	     �&  �	     �&  �	     )'   �	     T'  $�	     �'  (�	     �'  ,�	     �'  0�	     (  4�	     %(  8�	     <(  <�	     O(  @�	     a(  D�	     y(  H�	     �(  L�	     �(  P�	     �(  T�	     �(  X�	     �(  \�	     )  `�	     )  d�	     +)  h�	     D)  l�	     ])  p�	     p)  t�	     �)  x�	     �)  |�	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ċ	     �+  ȋ	     �+  ̋	     �+  Ћ	     ,  ԋ	     2,  ؋	     O,  ܋	     q,  ��	     �,  �	     �,  �	     �,  �	     �,  ��	     -  �	     --  ��	     Q-  ��	     t-   �	     �-  �	     �-  �	     �-  �	     .  �	     ,.  �	     S.  �	     {.  �	     �.   �	     �.  $�	     �.  (�	     '/  ,�	     G/  0�	     �7           ���#  8�	     �#  9�	     �#  :�	     �#  ;�	     $  <�	     2$  @�	     C$  D�	     T$  H�	     e$  L�	     |$  P�	     �$  T�	     �$  X�	     �$  \�	     �$  `�	     �$  d�	     %  h�	     L%  l�	     �%  p�	     �%  x�	     �%  |�	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  Č	     O(  Ȍ	     a(  ̌	     y(  Ќ	     �(  Ԍ	     �(  ،	     �(  ܌	     �(  ��	     �(  �	     )  �	     )  �	     +)  ��	     D)  �	     ])  ��	     p)  ��	     �)   �	     �)  �	     �)  �	     �)  �	     �)  �	     �)  �	     *  �	     +*  �	     D*   �	     X*  $�	     m*  (�	     �*  ,�	     �*  0�	     �*  4�	     �*  8�	     �*  <�	     +  @�	     9+  D�	     ^+  H�	     +  L�	     �+  P�	     �+  T�	     �+  X�	     ,  \�	     2,  `�	     O,  d�	     q,  h�	     �,  l�	     �,  p�	     �,  t�	     �,  x�	     -  |�	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     8           ���#  ލ	     �#  ߍ	     �#  ��	     �#  �	     $  �	     2$  �	     C$  �	     T$  �	     e$  ��	     |$  �	     �$  ��	     �$  ��	     �$   �	     �$  �	     �$  �	     %  �	     L%  �	     �%  �	     �%   �	     �%  $�	     �%  (�	     �%  ,�	     &  0�	     =&  4�	     i&  8�	     �&  <�	     �&  @�	     �&  D�	     �&  H�	     �&  L�	     )'  P�	     T'  T�	     �'  X�	     �'  \�	     �'  `�	     (  d�	     %(  h�	     <(  l�	     O(  p�	     a(  t�	     y(  x�	     �(  |�	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  Ď	     D*  Ȏ	     X*  ̎	     m*  Ў	     �*  Ԏ	     �*  ؎	     �*  ܎	     �*  ��	     �*  �	     +  �	     9+  �	     ^+  ��	     +  �	     �+  ��	     �+  ��	     �+   �	     ,  �	     2,  �	     O,  �	     q,  �	     �,  �	     �,  �	     �,  �	     �,   �	     -  $�	     --  (�	     Q-  ,�	     t-  0�	     �-  4�	     �-  8�	     �-  <�	     .  @�	     ,.  D�	     S.  H�	     {.  L�	     �.  P�	     �.  T�	     �.  X�	     '/  \�	     G/  `�	     8           ���#  l�	     �#  m�	     �#  n�	     �#  o�	     $  p�	     2$  t�	     C$  x�	     T$  |�	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ď	     i&  ȏ	     �&  ̏	     �&  Џ	     �&  ԏ	     �&  ؏	     �&  ܏	     )'  ��	     T'  �	     �'  �	     �'  �	     �'  ��	     (  �	     %(  ��	     <(  ��	     O(   �	     a(  �	     y(  �	     �(  �	     �(  �	     �(  �	     �(  �	     �(  �	     )   �	     )  $�	     +)  (�	     D)  ,�	     ])  0�	     p)  4�	     �)  8�	     �)  <�	     �)  @�	     �)  D�	     �)  H�	     �)  L�	     *  P�	     +*  T�	     D*  X�	     X*  \�	     m*  `�	     �*  d�	     �*  h�	     �*  l�	     �*  p�	     �*  t�	     +  x�	     9+  |�	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  Đ	     �-  Ȑ	     �-  ̐	     .  А	     ,.  Ԑ	     S.  ؐ	     {.  ܐ	     �.  ��	     �.  �	     �.  �	     '/  �	     G/  �	     8           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$   �	     C$  �	     T$  �	     e$  �	     |$  �	     �$  �	     �$  �	     �$  �	     �$   �	     �$  $�	     %  (�	     L%  ,�	     �%  0�	     �%  8�	     �%  <�	     �%  @�	     �%  D�	     &  H�	     =&  L�	     i&  P�	     �&  T�	     �&  X�	     �&  \�	     �&  `�	     �&  d�	     )'  h�	     T'  l�	     �'  p�	     �'  t�	     �'  x�	     (  |�	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  đ	     �)  ȑ	     �)  ̑	     �)  Б	     �)  ԑ	     *  ؑ	     +*  ܑ	     D*  ��	     X*  �	     m*  �	     �*  �	     �*  �	     �*  ��	     �*  ��	     �*  ��	     +   �	     9+  �	     ^+  �	     +  �	     �+  �	     �+  �	     �+  �	     ,  �	     2,   �	     O,  $�	     q,  (�	     �,  ,�	     �,  0�	     �,  4�	     �,  8�	     -  <�	     --  @�	     Q-  D�	     t-  H�	     �-  L�	     �-  P�	     �-  T�	     .  X�	     ,.  \�	     S.  `�	     {.  d�	     �.  h�	     �.  l�	     �.  p�	     '/  t�	     G/  x�	     -8           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  Ē	     �%  Ȓ	     �%  ̒	     &  В	     =&  Ԓ	     i&  ؒ	     �&  ܒ	     �&  ��	     �&  �	     �&  �	     �&  �	     )'  �	     T'  ��	     �'  ��	     �'  ��	     �'   �	     (  �	     %(  �	     <(  �	     O(  �	     a(  �	     y(  �	     �(  �	     �(   �	     �(  $�	     �(  (�	     �(  ,�	     )  0�	     )  4�	     +)  8�	     D)  <�	     ])  @�	     p)  D�	     �)  H�	     �)  L�	     �)  P�	     �)  T�	     �)  X�	     �)  \�	     *  `�	     +*  d�	     D*  h�	     X*  l�	     m*  p�	     �*  t�	     �*  x�	     �*  |�	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ē	     --  ȓ	     Q-  ̓	     t-  Г	     �-  ԓ	     �-  ؓ	     �-  ܓ	     .  ��	     ,.  �	     S.  �	     {.  �	     �.  �	     �.  ��	     �.  ��	     '/  ��	     G/   �	     B8           ���#  �	     �#  	�	     �#  
�	     �#  �	     $  �	     2$  �	     C$  �	     T$  �	     e$  �	     |$   �	     �$  $�	     �$  (�	     �$  ,�	     �$  0�	     �$  4�	     %  8�	     L%  <�	     �%  @�	     �%  H�	     �%  L�	     �%  P�	     �%  T�	     &  X�	     =&  \�	     i&  `�	     �&  d�	     �&  h�	     �&  l�	     �&  p�	     �&  t�	     )'  x�	     T'  |�	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  Ĕ	     ])  Ȕ	     p)  ̔	     �)  Д	     �)  Ԕ	     �)  ؔ	     �)  ܔ	     �)  ��	     �)  �	     *  �	     +*  �	     D*  �	     X*  ��	     m*  ��	     �*  ��	     �*   �	     �*  �	     �*  �	     �*  �	     +  �	     9+  �	     ^+  �	     +  �	     �+   �	     �+  $�	     �+  (�	     ,  ,�	     2,  0�	     O,  4�	     q,  8�	     �,  <�	     �,  @�	     �,  D�	     �,  H�	     -  L�	     --  P�	     Q-  T�	     t-  X�	     �-  \�	     �-  `�	     �-  d�	     .  h�	     ,.  l�	     S.  p�	     {.  t�	     �.  x�	     �.  |�	     �.  ��	     '/  ��	     G/  ��	     Y8           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ĕ	     �%  ȕ	     �%  Е	     �%  ԕ	     �%  ؕ	     �%  ܕ	     &  ��	     =&  �	     i&  �	     �&  �	     �&  �	     �&  ��	     �&  ��	     �&  ��	     )'   �	     T'  �	     �'  �	     �'  �	     �'  �	     (  �	     %(  �	     <(  �	     O(   �	     a(  $�	     y(  (�	     �(  ,�	     �(  0�	     �(  4�	     �(  8�	     �(  <�	     )  @�	     )  D�	     +)  H�	     D)  L�	     ])  P�	     p)  T�	     �)  X�	     �)  \�	     �)  `�	     �)  d�	     �)  h�	     �)  l�	     *  p�	     +*  t�	     D*  x�	     X*  |�	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  Ė	     �,  Ȗ	     �,  ̖	     �,  Ж	     -  Ԗ	     --  ؖ	     Q-  ܖ	     t-  ��	     �-  �	     �-  �	     �-  �	     .  �	     ,.  ��	     S.  ��	     {.  ��	     �.   �	     �.  �	     �.  �	     '/  �	     G/  �	     q8           ���#  �	     �#  �	     �#  �	     �#  �	     $  �	     2$   �	     C$  $�	     T$  (�	     e$  ,�	     |$  0�	     �$  4�	     �$  8�	     �$  <�	     �$  @�	     �$  D�	     %  H�	     L%  L�	     �%  P�	     �%  X�	     �%  \�	     �%  `�	     �%  d�	     &  h�	     =&  l�	     i&  p�	     �&  t�	     �&  x�	     �&  |�	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ė	     )  ȗ	     )  ̗	     +)  З	     D)  ԗ	     ])  ؗ	     p)  ܗ	     �)  ��	     �)  �	     �)  �	     �)  �	     �)  �	     �)  ��	     *  ��	     +*  ��	     D*   �	     X*  �	     m*  �	     �*  �	     �*  �	     �*  �	     �*  �	     �*  �	     +   �	     9+  $�	     ^+  (�	     +  ,�	     �+  0�	     �+  4�	     �+  8�	     ,  <�	     2,  @�	     O,  D�	     q,  H�	     �,  L�	     �,  P�	     �,  T�	     �,  X�	     -  \�	     --  `�	     Q-  d�	     t-  h�	     �-  l�	     �-  p�	     �-  t�	     .  x�	     ,.  |�	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �8           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  Ę	     �$  Ș	     �$  ̘	     %  И	     L%  Ԙ	     �%  ؘ	     �%  ��	     �%  �	     �%  �	     �%  �	     &  �	     =&  ��	     i&  ��	     �&  ��	     �&   �	     �&  �	     �&  �	     �&  �	     )'  �	     T'  �	     �'  �	     �'  �	     �'   �	     (  $�	     %(  (�	     <(  ,�	     O(  0�	     a(  4�	     y(  8�	     �(  <�	     �(  @�	     �(  D�	     �(  H�	     �(  L�	     )  P�	     )  T�	     +)  X�	     D)  \�	     ])  `�	     p)  d�	     �)  h�	     �)  l�	     �)  p�	     �)  t�	     �)  x�	     �)  |�	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ę	     2,  ș	     O,  ̙	     q,  Й	     �,  ԙ	     �,  ؙ	     �,  ܙ	     �,  ��	     -  �	     --  �	     Q-  �	     t-  �	     �-  ��	     �-  ��	     �-  ��	     .   �	     ,.  �	     S.  �	     {.  �	     �.  �	     �.  �	     �.  �	     '/  �	     G/   �	     �8           ���#  (�	     �#  )�	     �#  *�	     �#  +�	     $  ,�	     2$  0�	     C$  4�	     T$  8�	     e$  <�	     |$  @�	     �$  D�	     �$  H�	     �$  L�	     �$  P�	     �$  T�	     %  X�	     L%  \�	     �%  `�	     �%  h�	     �%  l�	     �%  p�	     �%  t�	     &  x�	     =&  |�	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  Ě	     �(  Ț	     �(  ̚	     �(  К	     �(  Ԛ	     )  ؚ	     )  ܚ	     +)  ��	     D)  �	     ])  �	     p)  �	     �)  �	     �)  ��	     �)  ��	     �)  ��	     �)   �	     �)  �	     *  �	     +*  �	     D*  �	     X*  �	     m*  �	     �*  �	     �*   �	     �*  $�	     �*  (�	     �*  ,�	     +  0�	     9+  4�	     ^+  8�	     +  <�	     �+  @�	     �+  D�	     �+  H�	     ,  L�	     2,  P�	     O,  T�	     q,  X�	     �,  \�	     �,  `�	     �,  d�	     �,  h�	     -  l�	     --  p�	     Q-  t�	     t-  x�	     �-  |�	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �8           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ě	     |$  ț	     �$  ̛	     �$  Л	     �$  ԛ	     �$  ؛	     �$  ܛ	     %  ��	     L%  �	     �%  �	     �%  �	     �%  ��	     �%  ��	     �%  ��	     &   �	     =&  �	     i&  �	     �&  �	     �&  �	     �&  �	     �&  �	     �&  �	     )'   �	     T'  $�	     �'  (�	     �'  ,�	     �'  0�	     (  4�	     %(  8�	     <(  <�	     O(  @�	     a(  D�	     y(  H�	     �(  L�	     �(  P�	     �(  T�	     �(  X�	     �(  \�	     )  `�	     )  d�	     +)  h�	     D)  l�	     ])  p�	     p)  t�	     �)  x�	     �)  |�	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  Ĝ	     �+  Ȝ	     �+  ̜	     �+  М	     ,  Ԝ	     2,  ؜	     O,  ܜ	     q,  ��	     �,  �	     �,  �	     �,  �	     �,  �	     -  ��	     --  ��	     Q-  ��	     t-   �	     �-  �	     �-  �	     �-  �	     .  �	     ,.  �	     S.  �	     {.  �	     �.   �	     �.  $�	     �.  (�	     '/  ,�	     G/  0�	     �8           ���#  8�	     �#  9�	     �#  :�	     �#  ;�	     $  <�	     2$  @�	     C$  D�	     T$  H�	     e$  L�	     |$  P�	     �$  T�	     �$  X�	     �$  \�	     �$  `�	     �$  d�	     %  h�	     L%  l�	     �%  p�	     �%  x�	     �%  |�	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ĝ	     O(  ȝ	     a(  ̝	     y(  Н	     �(  ԝ	     �(  ؝	     �(  ܝ	     �(  ��	     �(  �	     )  �	     )  �	     +)  �	     D)  ��	     ])  ��	     p)  ��	     �)   �	     �)  �	     �)  �	     �)  �	     �)  �	     �)  �	     *  �	     +*  �	     D*   �	     X*  $�	     m*  (�	     �*  ,�	     �*  0�	     �*  4�	     �*  8�	     �*  <�	     +  @�	     9+  D�	     ^+  H�	     +  L�	     �+  P�	     �+  T�	     �+  X�	     ,  \�	     2,  `�	     O,  d�	     q,  h�	     �,  l�	     �,  p�	     �,  t�	     �,  x�	     -  |�	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �8           ���#  ��	     �#  ��	     �#  	     �#  Þ	     $  Ğ	     2$  Ȟ	     C$  ̞	     T$  О	     e$  Ԟ	     |$  ؞	     �$  ܞ	     �$  ��	     �$  �	     �$  �	     �$  �	     %  �	     L%  ��	     �%  ��	     �%   �	     �%  �	     �%  �	     �%  �	     &  �	     =&  �	     i&  �	     �&  �	     �&   �	     �&  $�	     �&  (�	     �&  ,�	     )'  0�	     T'  4�	     �'  8�	     �'  <�	     �'  @�	     (  D�	     %(  H�	     <(  L�	     O(  P�	     a(  T�	     y(  X�	     �(  \�	     �(  `�	     �(  d�	     �(  h�	     �(  l�	     )  p�	     )  t�	     +)  x�	     D)  |�	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ğ	     +  ȟ	     9+  ̟	     ^+  П	     +  ԟ	     �+  ؟	     �+  ܟ	     �+  ��	     ,  �	     2,  �	     O,  �	     q,  �	     �,  ��	     �,  ��	     �,  ��	     �,   �	     -  �	     --  �	     Q-  �	     t-  �	     �-  �	     �-  �	     �-  �	     .   �	     ,.  $�	     S.  (�	     {.  ,�	     �.  0�	     �.  4�	     �.  8�	     '/  <�	     G/  @�	     �8           ���#  H�	     �#  I�	     �#  J�	     �#  K�	     $  L�	     2$  P�	     C$  T�	     T$  X�	     e$  \�	     |$  `�	     �$  d�	     �$  h�	     �$  l�	     �$  p�	     �$  t�	     %  x�	     L%  |�	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  Ġ	     �'  Ƞ	     (  ̠	     %(  Р	     <(  Ԡ	     O(  ؠ	     a(  ܠ	     y(  �	     �(  �	     �(  �	     �(  �	     �(  �	     �(  ��	     )  ��	     )  ��	     +)   �	     D)  �	     ])  �	     p)  �	     �)  �	     �)  �	     �)  �	     �)  �	     �)   �	     �)  $�	     *  (�	     +*  ,�	     D*  0�	     X*  4�	     m*  8�	     �*  <�	     �*  @�	     �*  D�	     �*  H�	     �*  L�	     +  P�	     9+  T�	     ^+  X�	     +  \�	     �+  `�	     �+  d�	     �+  h�	     ,  l�	     2,  p�	     O,  t�	     q,  x�	     �,  |�	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ġ	     G/  ȡ	     �8           ��9  ��      �#  С	     �#  ѡ	     �#  ҡ	     �#  ӡ	     $  ԡ	     2$  ء	     C$  ܡ	     T$  �	     e$  �	     |$  �	     �$  �	     �$  �	     �$  ��	     �$  ��	     �$  ��	     %   �	     L%  �	     �%  �	     �%  �	     �%  �	     �%  �	     �%  �	     &   �	     =&  $�	     i&  (�	     �&  ,�	     �&  0�	     �&  4�	     �&  8�	     �&  <�	     )'  @�	     T'  D�	     �'  H�	     �'  L�	     �'  P�	     (  T�	     %(  X�	     <(  \�	     O(  `�	     a(  d�	     y(  h�	     �(  l�	     �(  p�	     �(  t�	     �(  x�	     �(  |�	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  Ģ	     �*  Ȣ	     �*  ̢	     �*  Т	     �*  Ԣ	     +  آ	     9+  ܢ	     ^+  �	     +  �	     �+  �	     �+  �	     �+  �	     ,  ��	     2,  ��	     O,  ��	     q,   �	     �,  �	     �,  �	     �,  �	     �,  �	     -  �	     --  �	     Q-  �	     t-   �	     �-  $�	     �-  (�	     �-  ,�	     .  0�	     ,.  4�	     S.  8�	     {.  <�	     �.  @�	     �.  D�	     �.  H�	     '/  L�	     G/  P�	     99           ��G9  ��     �#  X�	     �#  Y�	     �#  Z�	     �#  [�	     $  \�	     2$  `�	     C$  d�	     T$  h�	     e$  l�	     |$  p�	     �$  t�	     �$  x�	     �$  |�	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ģ	     )'  ȣ	     T'  ̣	     �'  У	     �'  ԣ	     �'  أ	     (  ܣ	     %(  �	     <(  �	     O(  �	     a(  �	     y(  �	     �(  ��	     �(  ��	     �(  ��	     �(   �	     �(  �	     )  �	     )  �	     +)  �	     D)  �	     ])  �	     p)  �	     �)   �	     �)  $�	     �)  (�	     �)  ,�	     �)  0�	     �)  4�	     *  8�	     +*  <�	     D*  @�	     X*  D�	     m*  H�	     �*  L�	     �*  P�	     �*  T�	     �*  X�	     �*  \�	     +  `�	     9+  d�	     ^+  h�	     +  l�	     �+  p�	     �+  t�	     �+  x�	     ,  |�	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  Ĥ	     �.  Ȥ	     �.  ̤	     �.  Ф	     '/  Ԥ	     G/  ؤ	     o9           ���#  �	     �#  �	     �#  �	     �#  �	     $  �	     2$  �	     C$  �	     T$  �	     e$  ��	     |$  ��	     �$  ��	     �$   �	     �$  �	     �$  �	     �$  �	     %  �	     L%  �	     �%  �	     �%   �	     �%  $�	     �%  (�	     �%  ,�	     &  0�	     =&  4�	     i&  8�	     �&  <�	     �&  @�	     �&  D�	     �&  H�	     �&  L�	     )'  P�	     T'  T�	     �'  X�	     �'  \�	     �'  `�	     (  d�	     %(  h�	     <(  l�	     O(  p�	     a(  t�	     y(  x�	     �(  |�	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ĥ	     D*  ȥ	     X*  ̥	     m*  Х	     �*  ԥ	     �*  إ	     �*  ܥ	     �*  �	     �*  �	     +  �	     9+  �	     ^+  �	     +  ��	     �+  ��	     �+  ��	     �+   �	     ,  �	     2,  �	     O,  �	     q,  �	     �,  �	     �,  �	     �,  �	     �,   �	     -  $�	     --  (�	     Q-  ,�	     t-  0�	     �-  4�	     �-  8�	     �-  <�	     .  @�	     ,.  D�	     S.  H�	     {.  L�	     �.  P�	     �.  T�	     �.  X�	     '/  \�	     G/  `�	     |9           ���#  h�	     �#  i�	     �#  j�	     �#  k�	     $  l�	     2$  p�	     C$  t�	     T$  x�	     e$  |�	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  Ħ	     �&  Ȧ	     �&  ̦	     �&  Ц	     �&  Ԧ	     )'  ئ	     T'  ܦ	     �'  �	     �'  �	     �'  �	     (  �	     %(  �	     <(  ��	     O(  ��	     a(  ��	     y(   �	     �(  �	     �(  �	     �(  �	     �(  �	     �(  �	     )  �	     )  �	     +)   �	     D)  $�	     ])  (�	     p)  ,�	     �)  0�	     �)  4�	     �)  8�	     �)  <�	     �)  @�	     �)  D�	     *  H�	     +*  L�	     D*  P�	     X*  T�	     m*  X�	     �*  \�	     �*  `�	     �*  d�	     �*  h�	     �*  l�	     +  p�	     9+  t�	     ^+  x�	     +  |�	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ħ	     .  ȧ	     ,.  ̧	     S.  Ч	     {.  ԧ	     �.  ا	     �.  ܧ	     �.  �	     '/  �	     G/  �	     �9           ���#  �	     �#  �	     �#  �	     �#  �	     $  ��	     2$  ��	     C$  ��	     T$   �	     e$  �	     |$  �	     �$  �	     �$  �	     �$  �	     �$  �	     �$  �	     %   �	     L%  $�	     �%  (�	     �%  0�	     �%  4�	     �%  8�	     �%  <�	     &  @�	     =&  D�	     i&  H�	     �&  L�	     �&  P�	     �&  T�	     �&  X�	     �&  \�	     )'  `�	     T'  d�	     �'  h�	     �'  l�	     �'  p�	     (  t�	     %(  x�	     <(  |�	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  Ĩ	     �)  Ȩ	     �)  ̨	     *  Ш	     +*  Ԩ	     D*  ب	     X*  ܨ	     m*  �	     �*  �	     �*  �	     �*  �	     �*  �	     �*  ��	     +  ��	     9+  ��	     ^+   �	     +  �	     �+  �	     �+  �	     �+  �	     ,  �	     2,  �	     O,  �	     q,   �	     �,  $�	     �,  (�	     �,  ,�	     �,  0�	     -  4�	     --  8�	     Q-  <�	     t-  @�	     �-  D�	     �-  H�	     �-  L�	     .  P�	     ,.  T�	     S.  X�	     {.  \�	     �.  `�	     �.  d�	     �.  h�	     '/  l�	     G/  p�	     �9           ���#  x�	     �#  y�	     �#  z�	     �#  {�	     $  |�	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ĩ	     &  ȩ	     =&  ̩	     i&  Щ	     �&  ԩ	     �&  ة	     �&  ܩ	     �&  �	     �&  �	     )'  �	     T'  �	     �'  �	     �'  ��	     �'  ��	     (  ��	     %(   �	     <(  �	     O(  �	     a(  �	     y(  �	     �(  �	     �(  �	     �(  �	     �(   �	     �(  $�	     )  (�	     )  ,�	     +)  0�	     D)  4�	     ])  8�	     p)  <�	     �)  @�	     �)  D�	     �)  H�	     �)  L�	     �)  P�	     �)  T�	     *  X�	     +*  \�	     D*  `�	     X*  d�	     m*  h�	     �*  l�	     �*  p�	     �*  t�	     �*  x�	     �*  |�	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  Ī	     t-  Ȫ	     �-  ̪	     �-  Ъ	     �-  Ԫ	     .  ت	     ,.  ܪ	     S.  �	     {.  �	     �.  �	     �.  �	     �.  �	     '/  ��	     G/  ��	     �9           ���#  �	     �#  �	     �#   �	     �#  !�	     $  "�	     2$  $�	     C$  (�	     T$  ,�	     e$  0�	     |$  4�	     �$  8�	     �$  <�	     �$  @�	     �$  D�	     �$  H�	     %  L�	     L%  P�	     �%  X�	     �%  `�	     �%  d�	     �%  h�	     �%  l�	     &  p�	     =&  t�	     i&  x�	     �&  |�	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ī	     �(  ȫ	     �(  ̫	     )  Ы	     )  ԫ	     +)  ث	     D)  ܫ	     ])  �	     p)  �	     �)  �	     �)  �	     �)  �	     �)  ��	     �)  ��	     �)  ��	     *   �	     +*  �	     D*  �	     X*  �	     m*  �	     �*  �	     �*  �	     �*  �	     �*   �	     �*  $�	     +  (�	     9+  ,�	     ^+  0�	     +  4�	     �+  8�	     �+  <�	     �+  @�	     ,  D�	     2,  H�	     O,  L�	     q,  P�	     �,  T�	     �,  X�	     �,  \�	     �,  `�	     -  d�	     --  h�	     Q-  l�	     t-  p�	     �-  t�	     �-  x�	     �-  |�	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �9           ���#  Ƭ	     �#  Ǭ	     �#  Ȭ	     �#  ɬ	     $  ʬ	     2$  ̬	     C$  Ь	     T$  Ԭ	     e$  ج	     |$  ܬ	     �$  �	     �$  �	     �$  �	     �$  �	     �$  �	     %  ��	     L%  ��	     �%   �	     �%  �	     �%  �	     �%  �	     �%  �	     &  �	     =&  �	     i&   �	     �&  $�	     �&  (�	     �&  ,�	     �&  0�	     �&  4�	     )'  8�	     T'  <�	     �'  @�	     �'  D�	     �'  H�	     (  L�	     %(  P�	     <(  T�	     O(  X�	     a(  \�	     y(  `�	     �(  d�	     �(  h�	     �(  l�	     �(  p�	     �(  t�	     )  x�	     )  |�	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ĭ	     �*  ȭ	     �*  ̭	     +  Э	     9+  ԭ	     ^+  ح	     +  ܭ	     �+  �	     �+  �	     �+  �	     ,  �	     2,  �	     O,  ��	     q,  ��	     �,  ��	     �,   �	     �,  �	     �,  �	     -  �	     --  �	     Q-  �	     t-  �	     �-  �	     �-   �	     �-  $�	     .  (�	     ,.  ,�	     S.  0�	     {.  4�	     �.  8�	     �.  <�	     �.  @�	     '/  D�	     G/  H�	     �9           ���#  P�	     �#  Q�	     �#  R�	     �#  S�	     $  T�	     2$  X�	     C$  \�	     T$  `�	     e$  d�	     |$  h�	     �$  l�	     �$  p�	     �$  t�	     �$  x�	     �$  |�	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  Į	     �'  Ȯ	     �'  ̮	     �'  Ю	     (  Ԯ	     %(  خ	     <(  ܮ	     O(  �	     a(  �	     y(  �	     �(  �	     �(  �	     �(  ��	     �(  ��	     �(  ��	     )   �	     )  �	     +)  �	     D)  �	     ])  �	     p)  �	     �)  �	     �)  �	     �)   �	     �)  $�	     �)  (�	     �)  ,�	     *  0�	     +*  4�	     D*  8�	     X*  <�	     m*  @�	     �*  D�	     �*  H�	     �*  L�	     �*  P�	     �*  T�	     +  X�	     9+  \�	     ^+  `�	     +  d�	     �+  h�	     �+  l�	     �+  p�	     ,  t�	     2,  x�	     O,  |�	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  į	     �.  ȯ	     '/  ̯	     G/  Я	     �9           ���#  د	     �#  ٯ	     �#  گ	     �#  ۯ	     $  ܯ	     2$  �	     C$  �	     T$  �	     e$  �	     |$  �	     �$  ��	     �$  ��	     �$  ��	     �$   �	     �$  �	     %  �	     L%  �	     �%  �	     �%  �	     �%  �	     �%   �	     �%  $�	     &  (�	     =&  ,�	     i&  0�	     �&  4�	     �&  8�	     �&  <�	     �&  @�	     �&  D�	     )'  H�	     T'  L�	     �'  P�	     �'  T�	     �'  X�	     (  \�	     %(  `�	     <(  d�	     O(  h�	     a(  l�	     y(  p�	     �(  t�	     �(  x�	     �(  |�	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  İ	     m*  Ȱ	     �*  ̰	     �*  а	     �*  ԰	     �*  ذ	     �*  ܰ	     +  �	     9+  �	     ^+  �	     +  �	     �+  �	     �+  ��	     �+  ��	     ,  ��	     2,   �	     O,  �	     q,  �	     �,  �	     �,  �	     �,  �	     �,  �	     -  �	     --   �	     Q-  $�	     t-  (�	     �-  ,�	     �-  0�	     �-  4�	     .  8�	     ,.  <�	     S.  @�	     {.  D�	     �.  H�	     �.  L�	     �.  P�	     '/  T�	     G/  X�	     �9           ���#  `�	     �#  a�	     �#  b�	     �#  c�	     $  d�	     2$  h�	     C$  l�	     T$  p�	     e$  t�	     |$  x�	     �$  |�	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ı	     �&  ȱ	     �&  ̱	     )'  б	     T'  Ա	     �'  ر	     �'  ܱ	     �'  �	     (  �	     %(  �	     <(  �	     O(  �	     a(  ��	     y(  ��	     �(  ��	     �(   �	     �(  �	     �(  �	     �(  �	     )  �	     )  �	     +)  �	     D)  �	     ])   �	     p)  $�	     �)  (�	     �)  ,�	     �)  0�	     �)  4�	     �)  8�	     �)  <�	     *  @�	     +*  D�	     D*  H�	     X*  L�	     m*  P�	     �*  T�	     �*  X�	     �*  \�	     �*  `�	     �*  d�	     +  h�	     9+  l�	     ^+  p�	     +  t�	     �+  x�	     �+  |�	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  Ĳ	     S.  Ȳ	     {.  ̲	     �.  в	     �.  Բ	     �.  ز	     '/  ܲ	     G/  �	     �9           ���#  �	     �#  �	     �#  �	     �#  �	     $  �	     2$  �	     C$  ��	     T$  ��	     e$  ��	     |$   �	     �$  �	     �$  �	     �$  �	     �$  �	     �$  �	     %  �	     L%  �	     �%   �	     �%  (�	     �%  ,�	     �%  0�	     �%  4�	     &  8�	     =&  <�	     i&  @�	     �&  D�	     �&  H�	     �&  L�	     �&  P�	     �&  T�	     )'  X�	     T'  \�	     �'  `�	     �'  d�	     �'  h�	     (  l�	     %(  p�	     <(  t�	     O(  x�	     a(  |�	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ĳ	     *  ȳ	     +*  ̳	     D*  г	     X*  Գ	     m*  س	     �*  ܳ	     �*  �	     �*  �	     �*  �	     �*  �	     +  �	     9+  ��	     ^+  ��	     +  ��	     �+   �	     �+  �	     �+  �	     ,  �	     2,  �	     O,  �	     q,  �	     �,  �	     �,   �	     �,  $�	     �,  (�	     -  ,�	     --  0�	     Q-  4�	     t-  8�	     �-  <�	     �-  @�	     �-  D�	     .  H�	     ,.  L�	     S.  P�	     {.  T�	     �.  X�	     �.  \�	     �.  `�	     '/  d�	     G/  h�	     �9           ���#  p�	     �#  q�	     �#  r�	     �#  s�	     $  t�	     2$  x�	     C$  |�	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  Ĵ	     i&  ȴ	     �&  ̴	     �&  д	     �&  Դ	     �&  ش	     �&  ܴ	     )'  �	     T'  �	     �'  �	     �'  �	     �'  �	     (  ��	     %(  ��	     <(  ��	     O(   �	     a(  �	     y(  �	     �(  �	     �(  �	     �(  �	     �(  �	     �(  �	     )   �	     )  $�	     +)  (�	     D)  ,�	     ])  0�	     p)  4�	     �)  8�	     �)  <�	     �)  @�	     �)  D�	     �)  H�	     �)  L�	     *  P�	     +*  T�	     D*  X�	     X*  \�	     m*  `�	     �*  d�	     �*  h�	     �*  l�	     �*  p�	     �*  t�	     +  x�	     9+  |�	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ĵ	     �-  ȵ	     �-  ̵	     .  е	     ,.  Ե	     S.  ص	     {.  ܵ	     �.  �	     �.  �	     �.  �	     '/  �	     G/  �	     �9           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$   �	     C$  �	     T$  �	     e$  �	     |$  �	     �$  �	     �$  �	     �$  �	     �$   �	     �$  $�	     %  (�	     L%  ,�	     �%  0�	     �%  8�	     �%  <�	     �%  @�	     �%  D�	     &  H�	     =&  L�	     i&  P�	     �&  T�	     �&  X�	     �&  \�	     �&  `�	     �&  d�	     )'  h�	     T'  l�	     �'  p�	     �'  t�	     �'  x�	     (  |�	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  Ķ	     �)  ȶ	     �)  ̶	     �)  ж	     �)  Զ	     *  ض	     +*  ܶ	     D*  �	     X*  �	     m*  �	     �*  �	     �*  �	     �*  ��	     �*  ��	     �*  ��	     +   �	     9+  �	     ^+  �	     +  �	     �+  �	     �+  �	     �+  �	     ,  �	     2,   �	     O,  $�	     q,  (�	     �,  ,�	     �,  0�	     �,  4�	     �,  8�	     -  <�	     --  @�	     Q-  D�	     t-  H�	     �-  L�	     �-  P�	     �-  T�	     .  X�	     ,.  \�	     S.  `�	     {.  d�	     �.  h�	     �.  l�	     �.  p�	     '/  t�	     G/  x�	     �9           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ķ	     �$  ȷ	     %  ̷	     L%  з	     �%  ط	     �%  �	     �%  �	     �%  �	     �%  �	     &  �	     =&  ��	     i&  ��	     �&  ��	     �&   �	     �&  �	     �&  �	     �&  �	     )'  �	     T'  �	     �'  �	     �'  �	     �'   �	     (  $�	     %(  (�	     <(  ,�	     O(  0�	     a(  4�	     y(  8�	     �(  <�	     �(  @�	     �(  D�	     �(  H�	     �(  L�	     )  P�	     )  T�	     +)  X�	     D)  \�	     ])  `�	     p)  d�	     �)  h�	     �)  l�	     �)  p�	     �)  t�	     �)  x�	     �)  |�	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ĸ	     2,  ȸ	     O,  ̸	     q,  и	     �,  Ը	     �,  ظ	     �,  ܸ	     �,  �	     -  �	     --  �	     Q-  �	     t-  �	     �-  ��	     �-  ��	     �-  ��	     .   �	     ,.  �	     S.  �	     {.  �	     �.  �	     �.  �	     �.  �	     '/  �	     G/   �	     :           ��:           ���#  4�	     �#  5�	     �#  6�	     �#  7�	     $  8�	     2$  <�	     C$  @�	     T$  D�	     e$  H�	     |$  L�	     �$  P�	     �$  T�	     �$  X�	     �$  \�	     �$  `�	     %  d�	     L%  h�	     �%  p�	     �%  x�	     �%  |�	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  Ĺ	     O(  ȹ	     a(  ̹	     y(  й	     �(  Թ	     �(  ع	     �(  ܹ	     �(  �	     �(  �	     )  �	     )  �	     +)  �	     D)  ��	     ])  ��	     p)  ��	     �)   �	     �)  �	     �)  �	     �)  �	     �)  �	     �)  �	     *  �	     +*  �	     D*   �	     X*  $�	     m*  (�	     �*  ,�	     �*  0�	     �*  4�	     �*  8�	     �*  <�	     +  @�	     9+  D�	     ^+  H�	     +  L�	     �+  P�	     �+  T�	     �+  X�	     ,  \�	     2,  `�	     O,  d�	     q,  h�	     �,  l�	     �,  p�	     �,  t�	     �,  x�	     -  |�	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     :           ���#  ��	     �#  ��	     �#  º	     �#  ú	     $  ĺ	     2$  Ⱥ	     C$  ̺	     T$  к	     e$  Ժ	     |$  غ	     �$  ܺ	     �$  �	     �$  �	     �$  �	     �$  �	     %  �	     L%  ��	     �%  ��	     �%   �	     �%  �	     �%  �	     �%  �	     &  �	     =&  �	     i&  �	     �&  �	     �&   �	     �&  $�	     �&  (�	     �&  ,�	     )'  0�	     T'  4�	     �'  8�	     �'  <�	     �'  @�	     (  D�	     %(  H�	     <(  L�	     O(  P�	     a(  T�	     y(  X�	     �(  \�	     �(  `�	     �(  d�	     �(  h�	     �(  l�	     )  p�	     )  t�	     +)  x�	     D)  |�	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  Ļ	     +  Ȼ	     9+  ̻	     ^+  л	     +  Ի	     �+  ػ	     �+  ܻ	     �+  �	     ,  �	     2,  �	     O,  �	     q,  �	     �,  ��	     �,  ��	     �,  ��	     �,   �	     -  �	     --  �	     Q-  �	     t-  �	     �-  �	     �-  �	     �-  �	     .   �	     ,.  $�	     S.  (�	     {.  ,�	     �.  0�	     �.  4�	     �.  8�	     '/  <�	     G/  @�	     %:           ���#  H�	     �#  I�	     �#  J�	     �#  K�	     $  L�	     2$  P�	     C$  T�	     T$  X�	     e$  \�	     |$  `�	     �$  d�	     �$  h�	     �$  l�	     �$  p�	     �$  t�	     %  x�	     L%  |�	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ļ	     �'  ȼ	     (  ̼	     %(  м	     <(  Լ	     O(  ؼ	     a(  ܼ	     y(  �	     �(  �	     �(  �	     �(  �	     �(  �	     �(  ��	     )  ��	     )  ��	     +)   �	     D)  �	     ])  �	     p)  �	     �)  �	     �)  �	     �)  �	     �)  �	     �)   �	     �)  $�	     *  (�	     +*  ,�	     D*  0�	     X*  4�	     m*  8�	     �*  <�	     �*  @�	     �*  D�	     �*  H�	     �*  L�	     +  P�	     9+  T�	     ^+  X�	     +  \�	     �+  `�	     �+  d�	     �+  h�	     ,  l�	     2,  p�	     O,  t�	     q,  x�	     �,  |�	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  Ľ	     G/  Ƚ	     1:           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$   �	     T$  �	     e$  �	     |$  �	     �$  �	     �$  �	     �$  �	     �$  �	     �$   �	     %  $�	     L%  (�	     �%  0�	     �%  8�	     �%  <�	     �%  @�	     �%  D�	     &  H�	     =&  L�	     i&  P�	     �&  T�	     �&  X�	     �&  \�	     �&  `�	     �&  d�	     )'  h�	     T'  l�	     �'  p�	     �'  t�	     �'  x�	     (  |�	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ľ	     �)  Ⱦ	     �)  ̾	     �)  о	     �)  Ծ	     *  ؾ	     +*  ܾ	     D*  �	     X*  �	     m*  �	     �*  �	     �*  �	     �*  ��	     �*  ��	     �*  ��	     +   �	     9+  �	     ^+  �	     +  �	     �+  �	     �+  �	     �+  �	     ,  �	     2,   �	     O,  $�	     q,  (�	     �,  ,�	     �,  0�	     �,  4�	     �,  8�	     -  <�	     --  @�	     Q-  D�	     t-  H�	     �-  L�	     �-  P�	     �-  T�	     .  X�	     ,.  \�	     S.  `�	     {.  d�	     �.  h�	     �.  l�	     �.  p�	     '/  t�	     G/  x�	     ;:           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  Ŀ	     �$  ȿ	     �$  ̿	     �$  п	     �$  Կ	     %  ؿ	     L%  ܿ	     �%  �	     �%  �	     �%  �	     �%  �	     �%  ��	     &  ��	     =&  ��	     i&   �	     �&  �	     �&  �	     �&  �	     �&  �	     �&  �	     )'  �	     T'  �	     �'   �	     �'  $�	     �'  (�	     (  ,�	     %(  0�	     <(  4�	     O(  8�	     a(  <�	     y(  @�	     �(  D�	     �(  H�	     �(  L�	     �(  P�	     �(  T�	     )  X�	     )  \�	     +)  `�	     D)  d�	     ])  h�	     p)  l�	     �)  p�	     �)  t�	     �)  x�	     �)  |�	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-   �	     �-  �	     .  �	     ,.  �	     S.  �	     {.  �	     �.  �	     �.  �	     �.   �	     '/  $�	     G/  (�	     H:           ���#  0�	     �#  1�	     �#  2�	     �#  3�	     $  4�	     2$  8�	     C$  <�	     T$  @�	     e$  D�	     |$  H�	     �$  L�	     �$  P�	     �$  T�	     �$  X�	     �$  \�	     %  `�	     L%  d�	     �%  h�	     �%  p�	     �%  t�	     �%  x�	     �%  |�	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)   �	     �)  �	     �)  �	     �)  �	     *  �	     +*  �	     D*  �	     X*  �	     m*   �	     �*  $�	     �*  (�	     �*  ,�	     �*  0�	     �*  4�	     +  8�	     9+  <�	     ^+  @�	     +  D�	     �+  H�	     �+  L�	     �+  P�	     ,  T�	     2,  X�	     O,  \�	     q,  `�	     �,  d�	     �,  h�	     �,  l�	     �,  p�	     -  t�	     --  x�	     Q-  |�	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     Q:           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%   �	     �%  �	     &  �	     =&  �	     i&  �	     �&  �	     �&  �	     �&  �	     �&   �	     �&  $�	     )'  (�	     T'  ,�	     �'  0�	     �'  4�	     �'  8�	     (  <�	     %(  @�	     <(  D�	     O(  H�	     a(  L�	     y(  P�	     �(  T�	     �(  X�	     �(  \�	     �(  `�	     �(  d�	     )  h�	     )  l�	     +)  p�	     D)  t�	     ])  x�	     p)  |�	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --   �	     Q-  �	     t-  �	     �-  �	     �-  �	     �-  �	     .  �	     ,.  �	     S.   �	     {.  $�	     �.  (�	     �.  ,�	     �.  0�	     '/  4�	     G/  8�	     [:           ���#  @�	     �#  A�	     �#  B�	     �#  C�	     $  D�	     2$  H�	     C$  L�	     T$  P�	     e$  T�	     |$  X�	     �$  \�	     �$  `�	     �$  d�	     �$  h�	     �$  l�	     %  p�	     L%  t�	     �%  x�	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])   �	     p)  �	     �)  �	     �)  �	     �)  �	     �)  �	     �)  �	     �)  �	     *   �	     +*  $�	     D*  (�	     X*  ,�	     m*  0�	     �*  4�	     �*  8�	     �*  <�	     �*  @�	     �*  D�	     +  H�	     9+  L�	     ^+  P�	     +  T�	     �+  X�	     �+  \�	     �+  `�	     ,  d�	     2,  h�	     O,  l�	     q,  p�	     �,  t�	     �,  x�	     �,  |�	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     e:           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%   �	     �%  �	     �%  �	     �%  �	     �%  �	     &  �	     =&  �	     i&   �	     �&  $�	     �&  (�	     �&  ,�	     �&  0�	     �&  4�	     )'  8�	     T'  <�	     �'  @�	     �'  D�	     �'  H�	     (  L�	     %(  P�	     <(  T�	     O(  X�	     a(  \�	     y(  `�	     �(  d�	     �(  h�	     �(  l�	     �(  p�	     �(  t�	     )  x�	     )  |�	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,   �	     �,  �	     �,  �	     -  �	     --  �	     Q-  �	     t-  �	     �-  �	     �-   �	     �-  $�	     .  (�	     ,.  ,�	     S.  0�	     {.  4�	     �.  8�	     �.  <�	     �.  @�	     '/  D�	     G/  H�	     n:           ���#  P�	     �#  Q�	     �#  R�	     �#  S�	     $  T�	     2$  X�	     C$  \�	     T$  `�	     e$  d�	     |$  h�	     �$  l�	     �$  p�	     �$  t�	     �$  x�	     �$  |�	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )   �	     )  �	     +)  �	     D)  �	     ])  �	     p)  �	     �)  �	     �)  �	     �)   �	     �)  $�	     �)  (�	     �)  ,�	     *  0�	     +*  4�	     D*  8�	     X*  <�	     m*  @�	     �*  D�	     �*  H�	     �*  L�	     �*  P�	     �*  T�	     +  X�	     9+  \�	     ^+  `�	     +  d�	     �+  h�	     �+  l�	     �+  p�	     ,  t�	     2,  x�	     O,  |�	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     w:           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$   �	     �$  �	     %  �	     L%  �	     �%  �	     �%  �	     �%  �	     �%   �	     �%  $�	     &  (�	     =&  ,�	     i&  0�	     �&  4�	     �&  8�	     �&  <�	     �&  @�	     �&  D�	     )'  H�	     T'  L�	     �'  P�	     �'  T�	     �'  X�	     (  \�	     %(  `�	     <(  d�	     O(  h�	     a(  l�	     y(  p�	     �(  t�	     �(  x�	     �(  |�	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,   �	     O,  �	     q,  �	     �,  �	     �,  �	     �,  �	     �,  �	     -  �	     --   �	     Q-  $�	     t-  (�	     �-  ,�	     �-  0�	     �-  4�	     .  8�	     ,.  <�	     S.  @�	     {.  D�	     �.  H�	     �.  L�	     �.  P�	     '/  T�	     G/  X�	     �:           ���#  `�	     �#  a�	     �#  b�	     �#  c�	     $  d�	     2$  h�	     C$  l�	     T$  p�	     e$  t�	     |$  x�	     �$  |�	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(   �	     �(  �	     �(  �	     �(  �	     )  �	     )  �	     +)  �	     D)  �	     ])   �	     p)  $�	     �)  (�	     �)  ,�	     �)  0�	     �)  4�	     �)  8�	     �)  <�	     *  @�	     +*  D�	     D*  H�	     X*  L�	     m*  P�	     �*  T�	     �*  X�	     �*  \�	     �*  `�	     �*  d�	     +  h�	     9+  l�	     ^+  p�	     +  t�	     �+  x�	     �+  |�	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �:           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$   �	     �$  �	     �$  �	     �$  �	     �$  �	     �$  �	     %  �	     L%  �	     �%   �	     �%  (�	     �%  ,�	     �%  0�	     �%  4�	     &  8�	     =&  <�	     i&  @�	     �&  D�	     �&  H�	     �&  L�	     �&  P�	     �&  T�	     )'  X�	     T'  \�	     �'  `�	     �'  d�	     �'  h�	     (  l�	     %(  p�	     <(  t�	     O(  x�	     a(  |�	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+   �	     �+  �	     �+  �	     ,  �	     2,  �	     O,  �	     q,  �	     �,  �	     �,   �	     �,  $�	     �,  (�	     -  ,�	     --  0�	     Q-  4�	     t-  8�	     �-  <�	     �-  @�	     �-  D�	     .  H�	     ,.  L�	     S.  P�	     {.  T�	     �.  X�	     �.  \�	     �.  `�	     '/  d�	     G/  h�	     �:           ���:  @k     �#  p�	     �#  q�	     �#  r�	     �#  s�	     $  t�	     2$  x�	     C$  |�	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(   �	     a(  �	     y(  �	     �(  �	     �(  �	     �(  �	     �(  �	     �(  �	     )   �	     )  $�	     +)  (�	     D)  ,�	     ])  0�	     p)  4�	     �)  8�	     �)  <�	     �)  @�	     �)  D�	     �)  H�	     �)  L�	     *  P�	     +*  T�	     D*  X�	     X*  \�	     m*  `�	     �*  d�	     �*  h�	     �*  l�	     �*  p�	     �*  t�	     +  x�	     9+  |�	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �:           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$   �	     C$  �	     T$  �	     e$  �	     |$  �	     �$  �	     �$  �	     �$  �	     �$   �	     �$  $�	     %  (�	     L%  ,�	     �%  0�	     �%  8�	     �%  <�	     �%  @�	     �%  D�	     &  H�	     =&  L�	     i&  P�	     �&  T�	     �&  X�	     �&  \�	     �&  `�	     �&  d�	     )'  h�	     T'  l�	     �'  p�	     �'  t�	     �'  x�	     (  |�	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +   �	     9+  �	     ^+  �	     +  �	     �+  �	     �+  �	     �+  �	     ,  �	     2,   �	     O,  $�	     q,  (�	     �,  ,�	     �,  0�	     �,  4�	     �,  8�	     -  <�	     --  @�	     Q-  D�	     t-  H�	     �-  L�	     �-  P�	     �-  T�	     .  X�	     ,.  \�	     S.  `�	     {.  d�	     �.  h�	     �.  l�	     �.  p�	     '/  t�	     G/  x�	     �:           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'   �	     (  �	     %(  �	     <(  �	     O(  �	     a(  �	     y(  �	     �(  �	     �(   �	     �(  $�	     �(  (�	     �(  ,�	     )  0�	     )  4�	     +)  8�	     D)  <�	     ])  @�	     p)  D�	     �)  H�	     �)  L�	     �)  P�	     �)  T�	     �)  X�	     �)  \�	     *  `�	     +*  d�	     D*  h�	     X*  l�	     m*  p�	     �*  t�	     �*  x�	     �*  |�	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/   �	     �:           ���#  �	     �#  	�	     �#  
�	     �#  �	     $  �	     2$  �	     C$  �	     T$  �	     e$  �	     |$   �	     �$  $�	     �$  (�	     �$  ,�	     �$  0�	     �$  4�	     %  8�	     L%  <�	     �%  @�	     �%  H�	     �%  L�	     �%  P�	     �%  T�	     &  X�	     =&  \�	     i&  `�	     �&  d�	     �&  h�	     �&  l�	     �&  p�	     �&  t�	     )'  x�	     T'  |�	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*   �	     �*  �	     �*  �	     �*  �	     +  �	     9+  �	     ^+  �	     +  �	     �+   �	     �+  $�	     �+  (�	     ,  ,�	     2,  0�	     O,  4�	     q,  8�	     �,  <�	     �,  @�	     �,  D�	     �,  H�	     -  L�	     --  P�	     Q-  T�	     t-  X�	     �-  \�	     �-  `�	     �-  d�	     .  h�	     ,.  l�	     S.  p�	     {.  t�	     �.  x�	     �.  |�	     �.  ��	     '/  ��	     G/  ��	     �:           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'   �	     T'  �	     �'  �	     �'  �	     �'  �	     (  �	     %(  �	     <(  �	     O(   �	     a(  $�	     y(  (�	     �(  ,�	     �(  0�	     �(  4�	     �(  8�	     �(  <�	     )  @�	     )  D�	     +)  H�	     D)  L�	     ])  P�	     p)  T�	     �)  X�	     �)  \�	     �)  `�	     �)  d�	     �)  h�	     �)  l�	     *  p�	     +*  t�	     D*  x�	     X*  |�	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.   �	     �.  �	     �.  �	     '/  �	     G/  �	     ;           ���#  �	     �#  �	     �#  �	     �#  �	     $  �	     2$   �	     C$  $�	     T$  (�	     e$  ,�	     |$  0�	     �$  4�	     �$  8�	     �$  <�	     �$  @�	     �$  D�	     %  H�	     L%  L�	     �%  P�	     �%  X�	     �%  \�	     �%  `�	     �%  d�	     &  h�	     =&  l�	     i&  p�	     �&  t�	     �&  x�	     �&  |�	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*   �	     X*  �	     m*  �	     �*  �	     �*  �	     �*  �	     �*  �	     �*  �	     +   �	     9+  $�	     ^+  (�	     +  ,�	     �+  0�	     �+  4�	     �+  8�	     ,  <�	     2,  @�	     O,  D�	     q,  H�	     �,  L�	     �,  P�	     �,  T�	     �,  X�	     -  \�	     --  `�	     Q-  d�	     t-  h�	     �-  l�	     �-  p�	     �-  t�	     .  x�	     ,.  |�	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     ;           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&   �	     �&  �	     �&  �	     �&  �	     )'  �	     T'  �	     �'  �	     �'  �	     �'   �	     (  $�	     %(  (�	     <(  ,�	     O(  0�	     a(  4�	     y(  8�	     �(  <�	     �(  @�	     �(  D�	     �(  H�	     �(  L�	     )  P�	     )  T�	     +)  X�	     D)  \�	     ])  `�	     p)  d�	     �)  h�	     �)  l�	     �)  p�	     �)  t�	     �)  x�	     �)  |�	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .   �	     ,.  �	     S.  �	     {.  �	     �.  �	     �.  �	     �.  �	     '/  �	     G/   �	     ;           ��&;  ��[     ;;  =��     �#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$   �	     �$  �	     �$  �	     %  �	     L%  �	     �%  �	     �%   �	     �%  $�	     �%  (�	     �%  ,�	     &  0�	     =&  4�	     i&  8�	     �&  <�	     �&  @�	     �&  D�	     �&  H�	     �&  L�	     )'  P�	     T'  T�	     �'  X�	     �'  \�	     �'  `�	     (  d�	     %(  h�	     <(  l�	     O(  p�	     a(  t�	     y(  x�	     �(  |�	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+   �	     ,  �	     2,  �	     O,  �	     q,  �	     �,  �	     �,  �	     �,  �	     �,   �	     -  $�	     --  (�	     Q-  ,�	     t-  0�	     �-  4�	     �-  8�	     �-  <�	     .  @�	     ,.  D�	     S.  H�	     {.  L�	     �.  P�	     �.  T�	     �.  X�	     '/  \�	     G/  `�	     Z;           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'   �	     T'  �	     �'  �	     �'  �	     �'  �	     (  �	     %(  �	     <(  �	     O(   �	     a(  $�	     y(  (�	     �(  ,�	     �(  0�	     �(  4�	     �(  8�	     �(  <�	     )  @�	     )  D�	     +)  H�	     D)  L�	     ])  P�	     p)  T�	     �)  X�	     �)  \�	     �)  `�	     �)  d�	     �)  h�	     �)  l�	     *  p�	     +*  t�	     D*  x�	     X*  |�	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.   �	     �.  �	     �.  �	     '/  �	     G/  �	     f;           ��r;           ���#  �	     �#  �	     �#  �	     �#  �	     $  �	     2$   �	     C$  $�	     T$  (�	     e$  ,�	     |$  0�	     �$  4�	     �$  8�	     �$  <�	     �$  @�	     �$  D�	     %  H�	     L%  L�	     �%  P�	     �%  X�	     �%  \�	     �%  `�	     �%  d�	     &  h�	     =&  l�	     i&  p�	     �&  t�	     �&  x�	     �&  |�	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*   �	     X*  �	     m*  �	     �*  �	     �*  �	     �*  �	     �*  �	     �*  �	     +   �	     9+  $�	     ^+  (�	     +  ,�	     �+  0�	     �+  4�	     �+  8�	     ,  <�	     2,  @�	     O,  D�	     q,  H�	     �,  L�	     �,  P�	     �,  T�	     �,  X�	     -  \�	     --  `�	     Q-  d�	     t-  h�	     �-  l�	     �-  p�	     �-  t�	     .  x�	     ,.  |�	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �;           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&   �	     �&  �	     �&  �	     �&  �	     )'  �	     T'  �	     �'  �	     �'  �	     �'   �	     (  $�	     %(  (�	     <(  ,�	     O(  0�	     a(  4�	     y(  8�	     �(  <�	     �(  @�	     �(  D�	     �(  H�	     �(  L�	     )  P�	     )  T�	     +)  X�	     D)  \�	     ])  `�	     p)  d�	     �)  h�	     �)  l�	     �)  p�	     �)  t�	     �)  x�	     �)  |�	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .   �	     ,.  �	     S.  �	     {.  �	     �.  �	     �.  �	     �.  �	     '/  �	     G/   �	     �;           ���#  (�	     �#  )�	     �#  *�	     �#  +�	     $  ,�	     2$  0�	     C$  4�	     T$  8�	     e$  <�	     |$  @�	     �$  D�	     �$  H�	     �$  L�	     �$  P�	     �$  T�	     %  X�	     L%  \�	     �%  `�	     �%  h�	     �%  l�	     �%  p�	     �%  t�	     &  x�	     =&  |�	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)   �	     �)  �	     *  �	     +*  �	     D*  �	     X*  �	     m*  �	     �*  �	     �*   �	     �*  $�	     �*  (�	     �*  ,�	     +  0�	     9+  4�	     ^+  8�	     +  <�	     �+  @�	     �+  D�	     �+  H�	     ,  L�	     2,  P�	     O,  T�	     q,  X�	     �,  \�	     �,  `�	     �,  d�	     �,  h�	     -  l�	     --  p�	     Q-  t�	     t-  x�	     �-  |�	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �;           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &   �	     =&  �	     i&  �	     �&  �	     �&  �	     �&  �	     �&  �	     �&  �	     )'   �	     T'  $�	     �'  (�	     �'  ,�	     �'  0�	     (  4�	     %(  8�	     <(  <�	     O(  @�	     a(  D�	     y(  H�	     �(  L�	     �(  P�	     �(  T�	     �(  X�	     �(  \�	     )  `�	     )  d�	     +)  h�	     D)  l�	     ])  p�	     p)  t�	     �)  x�	     �)  |�	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-   �	     �-  �	     �-  �	     �-  �	     .  �	     ,.  �	     S.  �	     {.  �	     �.   �	     �.  $�	     �.  (�	     '/  ,�	     G/  0�	     �;           ���#  8�	     �#  9�	     �#  :�	     �#  ;�	     $  <�	     2$  @�	     C$  D�	     T$  H�	     e$  L�	     |$  P�	     �$  T�	     �$  X�	     �$  \�	     �$  `�	     �$  d�	     %  h�	     L%  l�	     �%  p�	     �%  x�	     �%  |�	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)   �	     �)  �	     �)  �	     �)  �	     �)  �	     �)  �	     *  �	     +*  �	     D*   �	     X*  $�	     m*  (�	     �*  ,�	     �*  0�	     �*  4�	     �*  8�	     �*  <�	     +  @�	     9+  D�	     ^+  H�	     +  L�	     �+  P�	     �+  T�	     �+  X�	     ,  \�	     2,  `�	     O,  d�	     q,  h�	     �,  l�	     �,  p�	     �,  t�	     �,  x�	     -  |�	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �;           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%   �	     �%  �	     �%  �	     �%  �	     &  �	     =&  �	     i&  �	     �&  �	     �&   �	     �&  $�	     �&  (�	     �&  ,�	     )'  0�	     T'  4�	     �'  8�	     �'  <�	     �'  @�	     (  D�	     %(  H�	     <(  L�	     O(  P�	     a(  T�	     y(  X�	     �(  \�	     �(  `�	     �(  d�	     �(  h�	     �(  l�	     )  p�	     )  t�	     +)  x�	     D)  |�	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,   �	     -  �	     --  �	     Q-  �	     t-  �	     �-  �	     �-  �	     �-  �	     .   �	     ,.  $�	     S.  (�	     {.  ,�	     �.  0�	     �.  4�	     �.  8�	     '/  <�	     G/  @�	     �;           ���#  H�	     �#  I�	     �#  J�	     �#  K�	     $  L�	     2$  P�	     C$  T�	     T$  X�	     e$  \�	     |$  `�	     �$  d�	     �$  h�	     �$  l�	     �$  p�	     �$  t�	     %  x�	     L%  |�	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)   �	     D)  �	     ])  �	     p)  �	     �)  �	     �)  �	     �)  �	     �)  �	     �)   �	     �)  $�	     *  (�	     +*  ,�	     D*  0�	     X*  4�	     m*  8�	     �*  <�	     �*  @�	     �*  D�	     �*  H�	     �*  L�	     +  P�	     9+  T�	     ^+  X�	     +  \�	     �+  `�	     �+  d�	     �+  h�	     ,  l�	     2,  p�	     O,  t�	     q,  x�	     �,  |�	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �;           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %   �	     L%  �	     �%  �	     �%  �	     �%  �	     �%  �	     �%  �	     &   �	     =&  $�	     i&  (�	     �&  ,�	     �&  0�	     �&  4�	     �&  8�	     �&  <�	     )'  @�	     T'  D�	     �'  H�	     �'  L�	     �'  P�	     (  T�	     %(  X�	     <(  \�	     O(  `�	     a(  d�	     y(  h�	     �(  l�	     �(  p�	     �(  t�	     �(  x�	     �(  |�	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,   �	     �,  �	     �,  �	     �,  �	     �,  �	     -  �	     --  �	     Q-  �	     t-   �	     �-  $�	     �-  (�	     �-  ,�	     .  0�	     ,.  4�	     S.  8�	     {.  <�	     �.  @�	     �.  D�	     �.  H�	     '/  L�	     G/  P�	     �;           ���#  X�	     �#  Y�	     �#  Z�	     �#  [�	     $  \�	     2$  `�	     C$  d�	     T$  h�	     e$  l�	     |$  p�	     �$  t�	     �$  x�	     �$  |�	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(   �	     �(  �	     )  �	     )  �	     +)  �	     D)  �	     ])  �	     p)  �	     �)   �	     �)  $�	     �)  (�	     �)  ,�	     �)  0�	     �)  4�	     *  8�	     +*  <�	     D*  @�	     X*  D�	     m*  H�	     �*  L�	     �*  P�	     �*  T�	     �*  X�	     �*  \�	     +  `�	     9+  d�	     ^+  h�	     +  l�	     �+  p�	     �+  t�	     �+  x�	     ,  |�	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     �;           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$   �	     �$  �	     �$  �	     �$  �	     %  �	     L%  �	     �%  �	     �%   �	     �%  $�	     �%  (�	     �%  ,�	     &  0�	     =&  4�	     i&  8�	     �&  <�	     �&  @�	     �&  D�	     �&  H�	     �&  L�	     )'  P�	     T'  T�	     �'  X�	     �'  \�	     �'  `�	     (  d�	     %(  h�	     <(  l�	     O(  p�	     a(  t�	     y(  x�	     �(  |�	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+   �	     ,  �	     2,  �	     O,  �	     q,  �	     �,  �	     �,  �	     �,  �	     �,   �	     -  $�	     --  (�	     Q-  ,�	     t-  0�	     �-  4�	     �-  8�	     �-  <�	     .  @�	     ,.  D�	     S.  H�	     {.  L�	     �.  P�	     �.  T�	     �.  X�	     '/  \�	     G/  `�	     <           ���#  h�	     �#  i�	     �#  j�	     �#  k�	     $  l�	     2$  p�	     C$  t�	     T$  x�	     e$  |�	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(   �	     �(  �	     �(  �	     �(  �	     �(  �	     �(  �	     )  �	     )  �	     +)   �	     D)  $�	     ])  (�	     p)  ,�	     �)  0�	     �)  4�	     �)  8�	     �)  <�	     �)  @�	     �)  D�	     *  H�	     +*  L�	     D*  P�	     X*  T�	     m*  X�	     �*  \�	     �*  `�	     �*  d�	     �*  h�	     �*  l�	     +  p�	     9+  t�	     ^+  x�	     +  |�	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     <           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$   �	     e$  �	     |$  �	     �$  �	     �$  �	     �$  �	     �$  �	     �$  �	     %   �	     L%  $�	     �%  (�	     �%  0�	     �%  4�	     �%  8�	     �%  <�	     &  @�	     =&  D�	     i&  H�	     �&  L�	     �&  P�	     �&  T�	     �&  X�	     �&  \�	     )'  `�	     T'  d�	     �'  h�	     �'  l�	     �'  p�	     (  t�	     %(  x�	     <(  |�	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+   �	     +  �	     �+  �	     �+  �	     �+  �	     ,  �	     2,  �	     O,  �	     q,   �	     �,  $�	     �,  (�	     �,  ,�	     �,  0�	     -  4�	     --  8�	     Q-  <�	     t-  @�	     �-  D�	     �-  H�	     �-  L�	     .  P�	     ,.  T�	     S.  X�	     {.  \�	     �.  `�	     �.  d�	     �.  h�	     '/  l�	     G/  p�	     <           ���#  x�	     �#  y�	     �#  z�	     �#  {�	     $  |�	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'  ��	     �'  ��	     �'  ��	     (  ��	     %(   �	     <(  �	     O(  �	     a(  �	     y(  �	     �(  �	     �(  �	     �(  �	     �(   �	     �(  $�	     )  (�	     )  ,�	     +)  0�	     D)  4�	     ])  8�	     p)  <�	     �)  @�	     �)  D�	     �)  H�	     �)  L�	     �)  P�	     �)  T�	     *  X�	     +*  \�	     D*  `�	     X*  d�	     m*  h�	     �*  l�	     �*  p�	     �*  t�	     �*  x�	     �*  |�	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.  ��	     '/  ��	     G/  ��	     !<           ���#   �	     �#  �	     �#  �	     �#  �	     $  �	     2$  �	     C$  �	     T$  �	     e$  �	     |$  �	     �$  �	     �$   �	     �$  $�	     �$  (�	     �$  ,�	     %  0�	     L%  4�	     �%  8�	     �%  @�	     �%  D�	     �%  H�	     �%  L�	     &  P�	     =&  T�	     i&  X�	     �&  \�	     �&  `�	     �&  d�	     �&  h�	     �&  l�	     )'  p�	     T'  t�	     �'  x�	     �'  |�	     �'  ��	     (  ��	     %(  ��	     <(  ��	     O(  ��	     a(  ��	     y(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     �(  ��	     )  ��	     )  ��	     +)  ��	     D)  ��	     ])  ��	     p)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     �)  ��	     *  ��	     +*  ��	     D*  ��	     X*  ��	     m*  ��	     �*  ��	     �*  ��	     �*  ��	     �*   �	     �*  �	     +  �	     9+  �	     ^+  �	     +  �	     �+  �	     �+  �	     �+   �	     ,  $�	     2,  (�	     O,  ,�	     q,  0�	     �,  4�	     �,  8�	     �,  <�	     �,  @�	     -  D�	     --  H�	     Q-  L�	     t-  P�	     �-  T�	     �-  X�	     �-  \�	     .  `�	     ,.  d�	     S.  h�	     {.  l�	     �.  p�	     �.  t�	     �.  x�	     '/  |�	     G/  ��	     +<           ���#  ��	     �#  ��	     �#  ��	     �#  ��	     $  ��	     2$  ��	     C$  ��	     T$  ��	     e$  ��	     |$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     �$  ��	     %  ��	     L%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     �%  ��	     &  ��	     =&  ��	     i&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     �&  ��	     )'  ��	     T'  ��	     �'   �	     �'  �	     �'  �	     (  �	     %(  �	     <(  �	     O(  �	     a(  �	     y(   �	     �(  $�	     �(  (�	     �(  ,�	     �(  0�	     �(  4�	     )  8�	     )  <�	     +)  @�	     D)  D�	     ])  H�	     p)  L�	     �)  P�	     �)  T�	     �)  X�	     �)  \�	     �)  `�	     �)  d�	     *  h�	     +*  l�	     D*  p�	     X*  t�	     m*  x�	     �*  |�	     �*  ��	     �*  ��	     �*  ��	     �*  ��	     +  ��	     9+  ��	     ^+  ��	     +  ��	     �+  ��	     �+  ��	     �+  ��	     ,  ��	     2,  ��	     O,  ��	     q,  ��	     �,  ��	     �,  ��	     �,  ��	     �,  ��	     -  ��	     --  ��	     Q-  ��	     t-  ��	     �-  ��	     �-  ��	     �-  ��	     .  ��	     ,.  ��	     S.  ��	     {.  ��	     �.  ��	     �.  ��	     �.   �	     '/  �	     G/  �	                  ��5<  <D      K<  �.     a<  ��B  "  r<  �@   "  }<  �	     �<  ��<     �<  �   "  �<  �    "  �<  0`
   "  &=  �   "  1=   	1   !  f=   ��    �=  ��     �=   �@   !   >  p�     >  �$     ->  (	   !  Y>  �T  "  �>  �#     �>  ��G   "  �>  @�   "  �>  `     �>  P�8   "  [?  �	2   !  �?  ��1     �?  P>J   "  �?   8   "  1@  ��     6@  �?   "  G@  `Q1   "  �@  y4�     �@  A	   !  �@   	(   ! �@  �   "  A  @^     #A  p-    4A  ͜J    EA  ��     jA  @�   "  �A  �	   !  �A  ��"   "  �A  �8   "  �A  �E   !  B  ��Z   "  ,B   @H   "  qB  p    �B  �
	   !  �B  �E     �B  ��R   "  C  �	   !  C  ��     ;C  `�m    JC  �   "  �C  �	<   !  �C     "  �C  @`
   "  �C  ���   "   D  H	   !  D  ��V     (D  �8   "  ]D  ��    !  ~D  �   "  �D  �GB     �D  ��     �D  ��   "  �D   E     E  �{   "  8E   �  "  XE  `��   "  �E  �1y     �E  0~6   "  F  �z   "  ?F   �"   "  TF  `    bF  `     �F  i\   "  �F  ��   "  �F  �     �F  ��   "   G  ���   "  G  �e  "  MG  02$   "  }G  ��0   "  �G  ��     �G  2   "  �G  �D     �G  0�   "  �G  �	   !  H  �     $H   �  "  2H  @�j   "  �H  0�   "  �H  ��`   "  I   ��     qI  �1   "  �I  �E     �I  P�8   "  J  ��     #J  F*    \J  �$     pJ  L	   !  �J  ��   "  �J  �
	   !  �J   ��     �J  �Qp   "  K  к   "  %K  0�>   "  BK  ,	   !  oK  `�I     �K  �$     �K  �   "  �K  0�   "  $L  p     @L  ��   "  RL  �8   "  �L  �*c    �L  ��     M  �	%   !  *M  @�(   !  1M  ��   !  KM  �-I   "  �M  h		     �M  )�8     �M  0 G   "  �M  �%    �M  �)      N  �T7   "  iN  $     �N  �   "  �N  �}6   "  �N  ��     �N  `�Q    KO  ��   "  �O  �		     �O  P�   "  �O   ��     P  ��l   "  rP  p�W  "  �P   �3   "  �P  p@p   "  'Q   �     AQ  @ L   "  vQ  &�Y     �Q   �   "  �Q  �	   !  �Q  ���   "  R  *�
     R  �  "  YR  ��    !  �R  ��m   "  �R  @�@   "  �R  �   "  �R  �   "  S  ��     *S   	(   ! dS  pS  "  �S  `�d   "  �S   `
   "  �S  ���   "  �S   �2   "  �S  вB     &T  �6c   "  [T  ���     cT  ��m   "  �T  �   "  �T  @	4   !  �T  ��   "  U  ��N   "  <U  �8   "  qU    	4   !  �U   �     �U   �    �U  �1     �U   �   !  �U  �	@   !  �U  p�   "  �U  p~6   "  >V  �	     WV  ��   !  �V  `
   "  �V  ��S   "  �V  �	   !  
W  l		     &W  	   !  6W  ��  "  OW  �|     ^W  p}6   "  sW  ��7   "  �W  ��!   "  �W  �L     �W  HE   !  X  0�   "  2X  �     @X  K/+     UX  ��Z   "  �X  �m     �X  		   !  �X  �B�  "  Y  P�   "  ]Y  �	   !  sY  p:   "  �Y  �)     �Y  P(     �Y  `�!   "  8Z  �!     RZ  � 	   !  eZ  �	   !  yZ  �/     �Z  0/     �Z  U�     �Z  09   "  �Z  �
	     �Z  ��    "  3[  p$     J[  @	(   !  �[  ��   !  �[  �	   !  �[  ��!   "  �[   0`     #\  `�;   !  b\  �E   !  �\  ��      �\  p�}   "  �\  @�   "  	]  �     #]  @�   !  E]  ��{    X]  ���   "  }]  �    �]  �	     �]  �		     �]  ���  "  @^  p     o^  a��     z^  :�-     �^  ���   "  �^  �H�   "  �^  �`  "  _  �     '_  ��   "  q_  ��-     v_  B	   !  �_  `�   "  �_  �	2   !  `  ���   "  `  ��c     `  P(     .`   $!     F`  �#   "  e`  -��     x`           ~`  P�2   "  �`  p�#     �`  ��      �`  Н�  "  aa  ��    "  sa  �)c    �a  �1   "  �a  (E     �a  l	     �a   �X   "  b  ��=   "  b  P=�   "  Gb  ��R   "  ab  ��   "  �b  ��>   "  	c  @y   "  @c  �9   "  |c  �R  "  �c  ��    �c  0�A     �c  �C     d  ��q   "  (d  d		     ?d  �	   !  ad   �     xd  ��g     �d  ��     �d  0)J     �d  H		     �d  ;�0     �d      "  �d  ��Z   "  �d  @�   "  *e  @�!     @e  :E   "  te  �     �e  ���   "  �e  ��>   "  �e  p�F   "  �e  ��   "  �e  @h     f  ��S   "  <f  ��H   "  df  ��!     wf  ��|   "  �f  `�   "  �f  �"R     �f  �"   "  g  `�  "  �g  �7   "  �g  ��   "  �g   	<   !   h  �	     h  �fX     "h   ��     8h  �8@   "  hh  ��&   "  �h   �   "  �h  �]�  "  i  p  "  ,i  ��     Di  �  "  `i  �	    !  gi   Y�     qi  ��   "  {i  P�L   "  �i  ��$   "  �i  �,     �i  P��    �i  ��   "  �i  �T
   "  2j  p     Jj  0�   "  Tj  ��      hj  `�d  "  �j   1     	k  /I   "  `k  ��H   "  �k  �0     �k  @�.  "  �k  ��'  "  �k  P�   "  l  �N�  "  ml  p	   !  �l  ��N   "  �l  �d�   "  �l  `�   "  m  ��5     m   Wo   "  im  �	   !  ~m  P��    �m  �    �m  ��     �m  j�B     �m  `�   "  �m  P   "  n  �	(   !  2n  �_
   "  gn  ��  "  �n  �k  "  �n  P   "  4o  І   "  To  `�m   "  to  ��  "  �o  �;     �o  ��m     �o  �D     �o  ��   !  �o   	   !  4p  P     `p  �    "  zp  `�   "  �p   �   "  �p  ��0   !  /q  � 	,   !  ]q  �.I   "  �q  �]     �q  �0      �q  0�:   "  ,r   �   "  Zr   	   !  nr  �   "  �r  P     �r  �D.     �r  �	(   ! s  �E   !  !s  ���     @s  �      Ss  �D8     ~s  4D    	 �s  PlV  "  �s  @�%   "  �s  �	�   !  t  �   !  t   G/   "  tt  �	   !  �t  ��     �t  @:     �t  @	(   !  �t  ��   "  6u  h	   !  `u  @�   "  �u   �u   "  �u  �Z  "  /v  0�   "  <v     "  Gv  P�   !  \v    	   !  sv  p��   "  �v  '3      �v  p�   "  w  �D.     .w  0�   !  Ow  @     iw  0@   "  �w  ��  "  �w  24     �w   S+   "  �w  `�   "  x  �.   "  3x  @   "  �x  �   "  �x  	   !  �x  0�'     �x  	   !  �x   }+   "  y  �	     1y  |�   !  Ky  ��   "  �y  �E   !  �y  ���   "  �y  P#�     #z  �   "  0z  �)     Pz  @C     �z  ;u    �z  �"	   !  �z  ��   "  �z  `>   "  �z  ���  "  �z  ���  "  {   9   "  B{  ��<   !  �{  P�i  "  �{  �	   !  �{  ��O   "  �{  Я�     |   �   "  |  �     |  �f�   "  _|   	,   !  ||  @'�    �|  H�?     �|  �@_  "  �|  �-�    }  0�   "  ,}  �     G}  p�>   "  \}  �)c    s}  @�   "  �}  ��a   "  �}  ��`     �}  L�   !  �}     "  �}   v   "  ?~  `9   "  s~  ��   "  �~   �j   "  �~  (	   !  �~  ��T     �~  )     �~  pE   !  .  @�
   "  <  ���  "  P  `��  "  e  @�G   "  �   ;   "  �  0�!   "  �   �   "  �  0D     �  \	     &�  Ч   "  a�  �+�    }�   ��     ��  `D     ��  0�!   "  ��  �h\   "  �  pD     !�  �t   "  c�  		   !  s�  �0!     ��  P�H   "  ��  ��     Ӂ  ?��     �   �E   "  �  ��z     G�  ��  "  V�  ��%     n�  �|   "  ��        ��   :     ��  ��&   "  �  p;   "  *�  K�  "  ��  g3;     ��  �	<   ! ��  ��L   "  Ճ  �g   "  �   �     ,�  �		     C�  ��   "  g�  ��s   "  u�  ��"   "  ��  3    ��  ��     Ȅ   �   !  τ  �Q     �   	    !  �  �	   !  >�  ��   "  ��  �	   !  ��  	       ��#     ۅ  Pc�   "  
�  P`K   "  S�  �V[   "  ��  0�    ��  T1     ��   2   "  ��  pi\   "  :�  0�   "  {�  `�   !  ��  ��      ��  �   "  ��  �E   !  �  ��   "  4�  ��!   "  w�  @�     ��  @�T   "  ��  @�   "  ��  k�D     ��  �%   "  ш  �	   !  �  ��   !  �  �38     �  ��I   "  B�  �%   "  S�  �]X     Z�  ��|   "     �%   "  ܉  �	   !  ��  �	'   !  �  ��}   "  .�  ��   "  L�  �	   !  ]�   I.   "  ��  �|
   "  ��  /�q     ��   )     ��  a�   !  ϊ  0	     �  �	(   ! ,�  p   "  j�  ��I    {�  0�  "  ��  ��8   "  �  ��4   "  Q�   V`    o�  �*L   "  Ɍ  �
	     ܌  �V`  "  �   L   "  K�  �"   "  v�   r=  "  ��  �+I   "  ,�  ���   "  >�  `�     W�  `�(   "  a�  `E   !  }�  �	<   !  ��  �1&     ��  *5     ˎ  ��J   "  �  (		   !  �  8	   !  �  Ё   "  �  `W(    @�  �@   "  ��  �    ˏ  ��   !  ޏ   	,   !  �  ��G   "  J�  @E   !  a�  �L   "  ��  0�   "  ɐ  @�@   "  Ӑ  �   "  �  ��     ��  P�u   �  Y��     �  �   !  �   �3   "  &�  ��*     9�  �:   "  b�  �	   !  v�   �a     Ǒ  ��W   "  �  ��     �  �J(  "  A�  p�     i�  ���   "  v�  `>   "  ��  �!     ��  �(L   "  ֒  5
	     ��  ж!     (�  �	     A�  P		     X�  �)     o�  ��   !  ��   ��   "  ��  ��   "  �  ���   "  )�  �
�   "  r�  ��a   "  ��  �9   ��  `2�   "  Ŕ  8	   !  ܔ  �   "  )�  �9     J�  Ь�     h�  E��    y�  �!	   !  ��  ��s   "  ��  �     ��  �c�   "  ו  �4#   "  �  P�   "  �  @	   !  C�  �/�  "  p�  0�   "  ��  �;   "  ږ  @�   "  �   	(   !  ��  `]�   "  5�  �#�     U�  p�  "  ��  p1   "  ��  �	     ח  ��   "  ��  �.%     �  @	(   ! 7�  ��     K�  ��|     [�  @�   "  ��  �	   !  ʘ  �38     Ә  �Q     ��  �   !  ��  `C     3�  0�     L�  ��      R�   E  "  ��  ��     ę  ��$   "  �  �!	   !   �  �V`    �  0=     /�  ��   "  Z�  ��   "  ��  @		     ��   $   "  Ӛ  ��!   "  �  �G   "  W�     "  ��  @3�   "  ś   �   "  �  p?�   "  �  ��A     :�  �R   "  r�  `�S   "  ��  p|   "  ��  ��!   "  Ҝ  0�S   "  �  �$�    ��  �     �  P�     (�  О   "  7�   ��    G�   �  "  `�   �   "  p�  ��     ��  �     ��  �D     ڝ  x 	   !  �  �{h   "  �  @��     ?�  @�!   "  P�  ��k  "  ��  ПH   "  ٞ  P�\   "  �  @�"   "  �  �)     B�  ��     L�  Ѐ   "  [�  �+V    r�  ��     ��  p"]     ��  �     ϟ  ��   "  �   Z   "  8�  ��     a�  @�   "  ��  @	�  "  �  P�%   "  ��  ��   "  <�  �     Z�  `��     s�  ��    ǡ  �0v     ��  @	"   !   �  ��*   !  N�  ��I     V�  �-I   "  ��  @�   "  ��  `		     ��  ���     ��  ��   !  ˢ  ���   "  ߢ  `1�   "  =�  � �  "  s�   ��    ��  �	   !  ��   [(  "  ڣ   �S   "  ��  5��      �  �    �  ��   "  @�  ��&   "  c�  �   "  q�  �g\   "  ��  ��   "  ɤ  ��   !  �  ��     ��  @�m   "  $�  0\(  "  e�  ��\     x�   *V    ��  �   !  ��  P�   "  ҥ  @�   "  �  ��   "  �  W�3     �   �    !  &�  @ �   "  ^�  `��   "  ��  pS  "  ��  �xX   "  �  `��     $�  @	(   !  Y�  ��     m�  ��     ��  �	   !  ��  ���     ��  ��$   "  �  �	   !  �  0�$   "  0�  �  "  L�  L   "  ��  �		     ��  @�:   !  ��  � 	   !  �  ��0   "  !�  ��     4�   �     H�   �!   !  m�  P     ��  ��  "  ��  �X�  "  ۩  P�F    ��  0  "  �  �  "  5�  ��<   "  ?�  ��#     E�  ~�)     M�  Њ   "  m�  d	   !  ��  0�S   "  ��  �     Ū  �.%     Ϊ  �    �  t		     �  �x[   "  N�  �     i�  �!   "  ��  ���   "  ��  �     �  Щ    "  ,�  �,I   "  W�  �5"   "  ��  ��   !  ��  �:   "  ֬  ��o   "  �   �X    V�  @"g     z�  �	   !  ��  �		     ��  �!     ƭ   )     �  ��     %�   X  "  ��  `     ��  �G     ͮ   �   "  �  0�   "  �  ��(   "  �   25   "  k�  0�   "  x�  �	   !  ��  P�   "  ��  i�  "  �  �/      ��   -    ��  �e   "  ��  ��     ϰ  p�2   "  %�  �E     8�  @{   "  o�  �b     {�  ��     ��  �     ̱  0�d   "  �  �9Z   "  �  �!     5�  �G     <�  ��'   "  H�  P76   "  |�  �L   "  ��  ��     ��  <   "  ²  @�    Ѳ  Щ    "  �  �|   "  ��  �	     �  �    ,�   	<   ! e�  lD     ��  �     ��  ��   "  ��  ��   "  г              �  �0!     ��  p��   "  �  0S1   "  T�  �   "  c�  �\�   "  ��  |�   !  ۴  p��   "  (�  Y�%     .�  ��     Y�  `^�  "  µ  �		     ۵  @�$   !  ��  `�&   "  /�  �E   !  Q�  ��&   "  z�  `1   "  ��  �  "  Ѷ   �s   "  �  �     "�  T		     6�  �   "  ^�   	@   !  �  $	   !  ��  0   "  ޷  `�X     �  �@   "  T�  P`K   "  ��   H^   "  Ҹ  �
	     �  �1   "  �  м�  "  ��  R�W     ��  @   "  ��  �	   !  �  ��   !  (�  �E   !  >�  �&   "  l�  P�`   "  ��  ��=     ��  ��  "  ��  L�e     �  �	   !  �   :   "  S�  P   "  �  �	     ��  �)     ��  ~�      ��  p�     ػ  `�    !  �  �		     0�  �D     6�  ��   !  M�  ��   !  g�   ,   "  ��  $�   !  ��  @a7   "  �  �%   "  ?�   <   "  k�  H�   !  ��  0�
   "  ��  p�   "  ɽ  |		     �  ��@   "  �   w=   "  �  $�     6�  ��   "  n�  ��7   "  پ   �   "  ��  ��   "  8�  `d;   "  ��       "  Ͽ  ��.   "  ܿ  ��   "  �  ��c     '�   "f     T�  ��&   "  ��   �(  "  ��  �	   !  ��  g�T     ��  0     ��  М+   "  ��   ��     ��  p�&   "  �  �    (�  p     @�  P+L   "  n�  �      u�  �54   "  ��  �	   !  ��  P�B     ��  0,�    ��   �   "  �  0   "   �  `�   "  -�  �	"   !  S�  0n     r�  �E   !  ��  `��   "  ��  �	   !  ��  �K  "  5�  ���   "  }�  �   "  ��  p�
   "  ��  �|   "  ��  P�B     ��  �.     ��  �     ��  ��     
�  @��   "  <�   	,   !  a�  ��     t�  ��   "  ��  d�   !  ��  ��6     ��  0}   "  ��  
�     ��  �	   !  ��   �   "  ��  PDD     �  ��   !  )�  m��     H�  ��,     O�  �   "  `�  ��     e�  ���   "  ��  ��K   "  ��  p��   "  ��  �r   "  �   8   "  {�   �X   "  ��  	�$    ��  ��   "  ��  �   "  ��  	   !  ��  tD     ��  ���     �  �"	   !  4�  �	   !  E�  k7  "  ��  x		     ��  P     ��  0   "  �  Ծ%     	�  p{     �  �3      $�  ��_     <�  ʴ      M�  �	   !  x�  ��   "  ��  ��8   "  ��  `�   "   �  P�&   "  N�  ��   "  ��  ��   "  ��   ��   "  ��  4q   "  ��  ��S   "  	�  �	(   ! �   �X   "  I�   �S   "  t�  Z�0     ��  ��   "  ��  XE   !  ��  @�   "  ��  �!	   !  ��  �E   !  �  @2  "  ��   �<     ��  @   "  ��   	(   ! ��  �_   "  )�  �     A�  +�]     I�  ��3   "  ]�  �4   "  ��  �C     ��  P   "  �  �]     �  ��"   "  )�  o��     6�  �	   !  ^�  �)!     ~�  ��  "  ��  ��   "  ��  �11     ��  @�#     ��  �b�   "  �  ��     �  �4d   "  q�  ��     ��  ��     ��  �		     ��  ��Q     @�  �B     Y�  0     u�  �   "  ��  P�%   "  ��  ���    ��  �
	   !  ��  @	&   !  ��  ���   "  ��  �}3   "  ��  @|   "  +�   �   !  M�  �+I   "  u�  �E   !  ��  ��4   "  ��  p�A   "  ��  hE   !  ;�  j4     H�  �   "  U�  @�!   "  ��  p�W     ��  P �    ��  l	   !  ��  �
  "  �   �<   !  X�   �I   "  ��  �	   !  ��  ��   "  ��  � �   "  �  @�!   "  �  �     :�  ��   !  M�  @�m   "  r�  �E   !  ��  �	   !  ��  ��  "  ��  �C     ��   �$   !  ��  �=b   "  �  ���   "  C�  |     Y�  @�&   "  {�  �S(  "  ��  P�!   "  �  $E     �  �1   "  w�  `��   "  ��  ��p     ��  ��   "  ��  C	   !  ��  P+6     ��  B�     �  �   "  V�  p	   !  }�  ��     ��  ��   !  ��  ��!     ��  �b     ��  ��     ��  ��     	�   ;   "  9�  ��B   "  P�  �E     h�  J�%     o�  0<!   "  ��  �1   "  ��  �A  "  0�  `     G�  0	   !  [�   c   r�  �>   "  ��  �2;     ��  �"    ��  p�>   "  #�  `�S   "  N�  �	   !  c�  ��     ��  
	   !  ��  ��  "  ��  �	     ��  �%   "  A�  ��    !  T�  `	   !  k�  P�   "  ��  �0;     ��  `:  "  M�  �@   "  ��  @�   "  ��   z   "  4�  ��%     L�  k�;     R�  �	   !  c�  ��     ��  p     ��  �		     ��  8		     ��  ��C   !  �  �)   "  T�  2   "  ��  �+W     ��  7�"     ��  ��     ��  p�   "  ��              �  ��@     �  ���     ;�  �4.     E�  �
	     Y�   ��     v�  �   "  ��  �	,   !  ��  p�c     ��  ��j   "  �  �    �  ��S   "  J�  pM  "  z�  ��M   "  ��   �  "  �  @GB     %�  ���	  "  ��  �	   !  ��  P�   "  ��  �;   "  ��  �   "  B�  �   "  ^�  �<|   "  ��  `	  "  ��  @��     ��  0�$   "  ��  �     ��  ��o     ��  ���     �  �D      #�  @GB     @�  0�   "  \�  P>J   "  ��  X		     ��  �.     ��   �   "  ��  `�  "  �   	(   !  K�  p$     b�  Ј[   "  x�  ?�2     �  �1   "  ��  0�#   "  ��  ��X     �  @   "  )�  >��    .�  	   !  D�   f  "  ��  p�>   "  ��  �w=   "  �  @Nr   "  Z�  0�   "  ��  p�   "  ��  `     	�  �   "  �  �     1�  9   "  k�  �		     �  �   !  ��  ��     ��   	)   !  ��  �	   !  �  `:   "  C�  	   !  V�  P9   "  ��  0�   "  ��  ��$   "  ��  ��     ��  H	   !  ��  Pza   "  .�  @	.   !  `�  ���   "  ��  `<p   "  ��  `�#     ��  ��     ��  [�*     �  �(�     (�  �v    2�  ��   "  >�  ��   "  z�  �     ��  @bX     ��  �	   !  ��  /     ��  ��#     ��  ��!     �  x	   !  )�  ��"     0�  @"	$   !  G�  �	   !  N�  P�`   "  ��  �
   "  ��  ��     ��  (	   !  ��  ��     ��  �GB     ��  m�     ��   �     ��  PG�   "  -�  @�S   "  R�  0�   "  p�   �9     w�  �(     ��  �s   "  ��  �   "  �  `�   "  F�  |�   !  ��  �     ��  �     ��  ���   "  ��  PyX   "  �  0�>   "  %�  p!     F�  �    "  `�  �)-     ��  �     ��  ��m   "  ��  ��   "  ��  �     ��  P�     �   �   "  &�  p�   "  6�  0+K    X�  �L   "  ��  `�%   "  ��  ��   "  �  �;   "  D�  `     a�  3      i�  p!     ��  �&T     ��  P�   !  ��  p�!   "  �  ��   "  -�  �	   !  F�  d	   !  l�  `'     ��  ��u    ��  x24     ��  PZ5   "  �  �dc   "  N�  �	(   ! ��  dD     ��  �	   !  ��  @�  "  ��  G3      ��  �8   "  r�  ��i   "  ��  0�     ��  �"	   !  ��  ���   "  ��  @	@   !  �  e�8     �  �   "  ,�  `L   "  a�  �a�   "  ��  P	   "  ��  P{_   "  ��  ��"   "  ��  `	    !  �  �:!   "  -�  Н   "  7�  p�"   "  b�  h"	   !  w�  �;   "  ��  P�  "  ��  К�   "  ��  �b   "  ��  q�c     ��  ��C   !  .�  U0;     A�  �~6   "  _�  e�   "  ��  ��6   "  ��  �		     �  ąE    �  @X�     #�   H    U�  �C     ��  ��   "  ��  �	   !  ��  �S    ��  ��P     �  �y�   "  @�   �P     ^�  @�  "  |�  ��   "  ��  @�   "  	�  `��     @�   .I   "  ��  �	     ��  @�7   "  ��  �a6   "  ��  P�L   "  �  �'*     D�  @X�   "  ��  ��     ��  0-2    ��  �     ��  �E   !  ��  ��
     ��  �      �  4	   !  9�  0#     L�  `��   "  m�  �T   "  ��  ��   "  ��  �    "  .�  ��!     X�  ��%   "  j�  `Dw   "  ��   �3   "  ��  0��  "  T�  P   "  ��  ��   !  ��  ��     ��  ޠV     ��  08B   "  ,�  �8     5�  �	   !  `�  !�)     h�  �Q   "  ��  �P     ��  0�   "  ��   ��   "  �   �S   "  "�  P�5   "  8�  0�l   "  x�  ��L   "  ��  �	4   !  ��  ` 	4   !  ��  �a�  "  9�  p	   !  M�  ��   "  ��  �P     ��  ��3     ��  ��!     ��  ��7   "  3  �   "  u  P+6     �  @	   !  �   �   "  �   �     �  ��"   "   @      �   !  d    "  � �(Y      0�   "  W -�@     o ��7   "  � ��#     � @�   "  � �!      o4
      �Z�     & ��:   !  d  �2   "  n ��#   "  x ��F   "  �      � ��6   !   �	,   !  0 �8   "  � @�E     � �
	     � �D     � p		     � ��N   "   p(L   "  a ��U     v @	   !  � @�V   "  � ��1     � �   "   �
	      p�   "  Q 4�   !  g �	   !  n :E   "  � p�W     � �L   "  �  �     � �   !  7 ��   !  T � 	   !  i �
  "  � 0-I   "  � ��F   "  � �L   "  - \		     E �D*    ~ @,I   "  � P�!   "  � ��     � ��_     � �|(   "  	 ��%   "  2	 D	     R	 ��N   "  t	 L		     �	 ��   "  �	 �V5   "  �	 �D    
 ��   "  F
 7�4     M
 P�   "  ]
 �/      m
 @	@   !  �
 �3     �
 ��   "  �
 P��   "    ��8      <�   !  F �	0   !  V �f     � �*     � ŵ+     � ���     � ��F   "  � ��   "  � �|   "  \ `	$   !  �  �   "  �  ��   "  � ���  "  � ��T   "  � 4�!     � ��   "  � �,I   "  B  �!   "  c �+�     @	@   !  � �   "  � ��"   "  � `(!      Y�5     & $     > ��     Z �    z ��   !  � �	     � �/!     � @�K   "   @!     ; �mV  "  } �E   !  �  @  "   ��?   "  O �	(   ! � �7N   "  � 8E     � �"R     �  �~     � ��   "  : p�   "  _ �E   !  � ��     � �
	     � `�      `   "   �;   "  Y  �S   "  � �!!     � o�   "  � � 
   "   �	   !  3 ��   "  e -�     l �i7  "  � ��:     � 	   !  � m  "  G �  "  c �!     � �c     � @�R   "  � �o�   "   ��#      p��  "  � @�S   "  � ���     � ��F     � p��   "  ! p�     :  	(   !  f `w=   "  � �D     � ��7     � ��m   "  � `��   "   P	   !  - @�   "  h @U8  "  � �
	     � �q�   "   �o    � ��"   "  � �L   "  � 0	   "  � �E      �   "  " T	     E 0�z     ^ �   "  �  �   "  � ;�;     � `�k  "  ?  N1   "  � 0�!     � �_   "  �  W`    � @_u   "  : ��m   "  _ �	   !  � pC     � �e   "  � �     � p�   "   �)     3 �   "  > @�$   "  H 0�   "  � l1+     � ��    � �a6   "  � �D      � `�   "  � 0E      P�     ( ��   "  S P�7   "  �  6�   "  � p	  "  Q �	   !  w P  "  � 4     � Hk      � |"	     �  �   "  � <		     �        p�   "  ) !E     ; �T`   "  � `��   "  � `	(   !  � )�  "  E  P5X   "  �  ��!   "  �  `   "  �  �0     ! p.I   "  A! ��   !  X!  �s   "  �! @   "  �! ���   "  �! �   "  �! �{   "  " ��   "  5"  �   "  E" ���
  "  �" ��   "  �" ��     # �7?   "  8# ��:  "  K# ��   "  ]# p@   "  �# ��     $ ���   "  t$ @�    �$  �     �$ ��Z   "  % p@p   "  \% @�K   "  �% �	   !  �% �Y�     �% ��S   "  �% P;   "  &  P�  "  T& Е   "  t& @�H   "  �& �
	     �& p>   "  '  ��   "  ' �E     8' 	   !  d' p��   "  �' p�v   "  �' Шz   "  �' ��"     �' 1�     ( �k    ( �		     %( p�   "  2( �	1   !  g( xE   !  ( P$o    �( 0�7   "  ) �W�  "  l) �	   !  �) ,E     �) �(     �) `/I   "  �) @8   "  R* p9   "  �* �>   "  �*       �* �?     �*  �_   "  �* ��$   "  + ��I   "  4+ k�-     9+ �	(   !  o+ `�   "  �+ $     �+ H	   !  �+ ��     , �y   "  J, �!~     {, ��:    �, ��   "  K- �D4  "  �- p�   !  �- (	     �- �	   !  �- p�   "  . p�   !  6. ��     N. �;   "  {. `�6   "  �. @9   "  �. ��   "  / �	   !  )/ �   "  v/ ��   !  �/ PDD     �/ �Q   "  �/ @1     �/ �2      0 P�   "  &0  �     H0  �"   "  q0 ��  "  �0 D		     �0 �Kb  "  �0 �>   "  �0 ��   "  '1 p�|   "  �1 �	(   !  �1 �j    �1  !     �1 ��   "  2 �:   "  ?2 ���   "  q2 ��
     x2 p   "  �2 ��   "  �2 �CJ     �2 �E   !  �2 �E   !  
3 ��K   "  E3 ��   "  �3  ��     �3 �za   "  4 �	     /4  �P     M4 @�    !  g4 ;2   "  �4 @g     �4  Z   "  �4 �   "  �4 `��     5  �
   "  S5 �E     s5 p�Z   "  �5 ��=   "  �5 ��<   !  �5  H     6 ��R   "  26 �@   "  p6 hD     �6  H  "  7 �  "  7 �X    (7 ��     :7 Ph\   "  7 �6     �7 �8   "  �7 �D     �7 0�K   "  �7 p  "  A8 p�!   "  M8 `�   "  r8 ���  "  �8 �	   !  9 4�'     9    "  [9 `��     |9 �	   !  �9 t��     �9 ��   "  �9 Њ   "  �9 1=     �9 N4     �9  x[   "  : �E   !  S: @  "  �: `�   "  �: �	   !  ; 	   !  ; ���	  "  �;  	(   ! �; �W(    �; �	   !  �; P�8   "  d< P�
   "  t< ��   "  �< ��     �< �~6   "  �< �     = �     = ��     8= `	'   !  c=  �%   "  m= ��4     �= ��     �= ���   "  �= �#     �= `�     > ��&   "  *> �	(   !  U> �	   !  i>     "  �>  �;   !  �> P�w   "  �> `��   "  ? ��g     !? 0�K   "  9?  �   "  �? �	   !  �? D	   !  �? ��     �? ��m   "  @ 0�     @ @	#   !  D@ �	     `@ ��     |@ *�A     �@ PB   "  �@     �@  `   "  A ��%   "  MA ٟ#     bA �E     �A `�    �A ��q  "  �A �_
   "  �A �:   "  B PE   !  SB v/"     WB �%   "  �B 0o�  "  C P|   "  8C P�   "  HC `�   "  ZC ��T     `C �$     {C             �C ��P     �C  (L   "  D \�   !  &D  �   "  dD 0�     zD v�J    �D `�|   "  �D P�   "  <E �>�   "  ~E �$     �E `��     �E  �   "  �E ��   "  F 0��   "  .F ��   "  =F  �   "  XF ��   "  �F @�7   "  �F  �s   "  �F �p�   "  *G P��     WG `�   "  pG �     |G ��k  "  �G @�   "  �G p�A   "  �G 0�3   "  �G �W(    �G ���   "  H 0   "  )H p{     <H �+K    XH �Zo   "  �H �CJ     �H O��     �H ,�   !  �H  �   "  I Rr   "  aI �		     wI �>   "  �I �	   !  �I ��     �I ��I     �I O��     �I `*W    J ��   "  %J �    "  aJ ��J   "  wJ 
�     �J p�   "  �J P}   "  �J _�      �J 0IN  "  �J  �   !  K  �Y     K p�9   "  ,K ��>   "  BK ���   "  iK  ��   "  �K �.   "  �K ��    "  �K �!	   !  �K ��  "  L �w=   "  2L  �&   "  `L ��   !  sL ��   "  �L ��   !  M ���     M Ю�  "  �M  	    !  �M @:     �M  +L   "  #N `��     ?N �   "  JN P   "  TN a�;     ]N �I     �N �	   !  �N �$    �N p�     �N  <   "  *O �8@   "  ZO �	   !  aO �     �O Y{�    �O  3?   "  �O �r    �O  �|   "  NP �     iP ��!     �P  
   "  �P ߧK    �P ��
     �P ��0  "  �P P��   "  Q  :     -Q �g\   "  sQ ��T   "   crtstuff.c THREAD_TYPE_MAIN THREAD_TYPE_SUB THREAD_TYPE_VM86 THREAD_PRIORITY_NORMAL THREAD_PRIORITY_IDLE FS_SEEK_SET FS_SEEK_CUR FS_SEEK_END FS_NODE_TYPE_NONE FS_NODE_TYPE_ROOT FS_NODE_TYPE_MOUNTPOINT FS_NODE_TYPE_FOLDER FS_NODE_TYPE_FILE FS_NODE_TYPE_PIPE FS_REGISTER_AS_DELEGATE_SUCCESSFUL FS_REGISTER_AS_DELEGATE_FAILED_EXISTING FS_REGISTER_AS_DELEGATE_FAILED_DELEGATE_CREATION FS_TRANSACTION_NO_REPEAT_ID FS_TRANSACTION_WAITING FS_TRANSACTION_FINISHED FS_TRANSACTION_REPEAT FS_CREATE_NODE_STATUS_CREATED FS_CREATE_NODE_STATUS_UPDATED FS_CREATE_NODE_STATUS_FAILED_NO_PARENT FS_DISCOVERY_SUCCESSFUL FS_DISCOVERY_NOT_FOUND FS_DISCOVERY_BUSY FS_DISCOVERY_ERROR FS_TASKED_DELEGATE_REQUEST_TYPE_DISCOVER FS_TASKED_DELEGATE_REQUEST_TYPE_READ FS_TASKED_DELEGATE_REQUEST_TYPE_WRITE FS_TASKED_DELEGATE_REQUEST_TYPE_GET_LENGTH FS_TASKED_DELEGATE_REQUEST_TYPE_READ_DIRECTORY FS_TASKED_DELEGATE_REQUEST_TYPE_OPEN FS_TASKED_DELEGATE_REQUEST_TYPE_CLOSE FS_OPEN_SUCCESSFUL FS_OPEN_NOT_FOUND FS_OPEN_ERROR FS_OPEN_BUSY FS_READ_SUCCESSFUL FS_READ_INVALID_FD FS_READ_BUSY FS_READ_ERROR FS_WRITE_SUCCESSFUL FS_WRITE_INVALID_FD FS_WRITE_NOT_SUPPORTED FS_WRITE_BUSY FS_WRITE_ERROR FS_CLOSE_SUCCESSFUL FS_CLOSE_INVALID_FD FS_CLOSE_BUSY FS_CLOSE_ERROR FS_SEEK_SUCCESSFUL FS_SEEK_INVALID_FD FS_SEEK_ERROR FS_TELL_SUCCESSFUL FS_TELL_INVALID_FD FS_LENGTH_SUCCESSFUL FS_LENGTH_INVALID_FD FS_LENGTH_NOT_FOUND FS_LENGTH_BUSY FS_LENGTH_ERROR FS_CLONEFD_SUCCESSFUL FS_CLONEFD_INVALID_SOURCE_FD FS_CLONEFD_ERROR FS_PIPE_SUCCESSFUL FS_PIPE_ERROR SET_WORKING_DIRECTORY_SUCCESSFUL SET_WORKING_DIRECTORY_NOT_A_FOLDER SET_WORKING_DIRECTORY_NOT_FOUND SET_WORKING_DIRECTORY_ERROR GET_WORKING_DIRECTORY_SUCCESSFUL GET_WORKING_DIRECTORY_SIZE_EXCEEDED GET_WORKING_DIRECTORY_ERROR FS_OPEN_DIRECTORY_SUCCESSFUL FS_OPEN_DIRECTORY_NOT_FOUND FS_OPEN_DIRECTORY_ERROR FS_READ_DIRECTORY_SUCCESSFUL FS_READ_DIRECTORY_EOD FS_READ_DIRECTORY_ERROR FS_DIRECTORY_REFRESH_SUCCESSFUL FS_DIRECTORY_REFRESH_ERROR FS_DIRECTORY_REFRESH_BUSY MESSAGE_SEND_MODE_BLOCKING MESSAGE_SEND_MODE_NON_BLOCKING MESSAGE_RECEIVE_MODE_BLOCKING MESSAGE_RECEIVE_MODE_NON_BLOCKING MESSAGE_SEND_STATUS_SUCCESSFUL MESSAGE_SEND_STATUS_QUEUE_FULL MESSAGE_SEND_STATUS_FAILED MESSAGE_SEND_STATUS_EXCEEDS_MAXIMUM MESSAGE_RECEIVE_STATUS_SUCCESSFUL MESSAGE_RECEIVE_STATUS_QUEUE_EMPTY MESSAGE_RECEIVE_STATUS_FAILED MESSAGE_RECEIVE_STATUS_FAILED_NOT_PERMITTED MESSAGE_RECEIVE_STATUS_EXCEEDS_BUFFER_SIZE MESSAGE_RECEIVE_STATUS_INTERRUPTED KERNQUERY_STATUS_SUCCESSFUL KERNQUERY_STATUS_UNKNOWN_ID __CTOR_LIST__ __DTOR_LIST__ __EH_FRAME_BEGIN__ __JCR_LIST__ deregister_tm_clones register_tm_clones __do_global_dtors_aux completed.5140 dtor_idx.5142 frame_dummy object.5152 __CTOR_END__ __FRAME_END__ __JCR_END__ __do_global_ctors_aux del_op.cc eh_personality.cc _ZL12read_sleb128PKhPl _ZL16get_adjusted_ptrPKSt9type_infoS1_PPv _ZL28read_encoded_value_with_basehjPKhPj _ZL15get_ttype_entryP16lsda_header_infom _ZL20check_exception_specP16lsda_header_infoPKSt9type_infoPvl _ZL21base_of_encoded_valuehP15_Unwind_Context _ZL17parse_lsda_headerP15_Unwind_ContextPKhP16lsda_header_info new_opv.cc eh_throw.cc _ZL23__gxx_exception_cleanup19_Unwind_Reason_CodeP17_Unwind_Exception eh_call.cc ostream-inst.cc misc-inst.cc istream.cc locale-inst.cc _ZNSs4_Rep10_M_disposeERKSaIcE.part.10 _ZNKSt5ctypeIcE5widenEc.part.25 _GLOBAL__sub_I_locale_inst.cc allocator-inst.cc ctype.cc ios_init.cc _ZNSt8ios_base4InitC2Ev.part.4 ext-inst.cc streambuf.cc sstream-inst.cc _ZNSs4_Rep10_M_disposeERKSaIcE.part.11 ios.cc _ZZNSt8ios_base6xallocEvE6_S_top locale_facets.cc locale.cc _ZGVZN12_GLOBAL__N_122get_locale_cache_mutexEvE18locale_cache_mutex streambuf-inst.cc ios-inst.cc codecvt.cc monetary_members.cc fstream-inst.cc string-inst.cc _ZNSs4_Rep10_M_disposeERKSaIcE.part.12 functexcept.cc _ZNSs4_Rep10_M_disposeERKSaIcE.part.0 regex.cc compatibility.cc bad_cast.cc vmi_class_type_info.cc del_opv.cc eh_globals.cc _ZL10eh_globals eh_catch.cc eh_exception.cc tinfo.cc class_type_info.cc bad_alloc.cc eh_terminate.cc guard.cc eh_alloc.cc _ZL14emergency_used _ZL16emergency_buffer _ZL15dependents_used _ZL17dependents_buffer new_op.cc bad_typeid.cc guard_error.cc pure.cc dyncast.cc eh_aux_runtime.cc si_class_type_info.cc vterminate.cc _ZZN9__gnu_cxx27__verbose_terminate_handlerEvE11terminating eh_type.cc bad_array_length.cc locale_init.cc _ZN12_GLOBAL__N_116get_locale_mutexEv.part.4 _ZGVZN12_GLOBAL__N_116get_locale_mutexEvE12locale_mutex _ZN12_GLOBAL__N_19cache_vecE _ZN12_GLOBAL__N_19facet_vecE _ZN12_GLOBAL__N_18name_vecE _ZN12_GLOBAL__N_16name_cE _ZN12_GLOBAL__N_17ctype_cE _ZN12_GLOBAL__N_19codecvt_cE _ZN12_GLOBAL__N_110numpunct_cE _ZN12_GLOBAL__N_116numpunct_cache_cE _ZN12_GLOBAL__N_19num_get_cE _ZN12_GLOBAL__N_19num_put_cE _ZN12_GLOBAL__N_19collate_cE _ZN12_GLOBAL__N_119moneypunct_cache_cfE _ZN12_GLOBAL__N_113moneypunct_cfE _ZN12_GLOBAL__N_119moneypunct_cache_ctE _ZN12_GLOBAL__N_113moneypunct_ctE _ZN12_GLOBAL__N_111money_get_cE _ZN12_GLOBAL__N_111money_put_cE _ZN12_GLOBAL__N_117timepunct_cache_cE _ZN12_GLOBAL__N_111timepunct_cE _ZN12_GLOBAL__N_110time_get_cE _ZN12_GLOBAL__N_110time_put_cE _ZN12_GLOBAL__N_110messages_cE _ZN12_GLOBAL__N_113c_locale_implE _ZNSt6locale13_S_initializeEv.part.7 _ZN12_GLOBAL__N_18c_localeE ios_failure.cc ctype_configure_char.cc collate_members.cc iostream-inst.cc numeric_members.cc istream-inst.cc ios_locale.cc basic_file.cc _ZN12_GLOBAL__N_1L6xwriteEiPKcl CSWTCH.15 messages_members.cc stdexcept.cc c++locale.cc _ZN9__gnu_cxxL14category_namesE time_members.cc functional.cc snprintf_lite.cc future.cc _ZNK12_GLOBAL__N_121future_error_category4nameEv _ZN12_GLOBAL__N_121future_error_categoryD2Ev _ZTVN12_GLOBAL__N_121future_error_categoryE _ZN12_GLOBAL__N_121future_error_categoryD1Ev _ZN12_GLOBAL__N_121future_error_categoryD0Ev _ZNK12_GLOBAL__N_121future_error_category7messageEi _ZGVZN12_GLOBAL__N_126__future_category_instanceEvE5__fec _ZZN12_GLOBAL__N_126__future_category_instanceEvE5__fec _ZTSN12_GLOBAL__N_121future_error_categoryE _ZTIN12_GLOBAL__N_121future_error_categoryE system_error.cc _ZNK12_GLOBAL__N_122generic_error_category4nameEv _ZNK12_GLOBAL__N_121system_error_category4nameEv _ZN12_GLOBAL__N_121system_error_categoryD2Ev _ZN12_GLOBAL__N_121system_error_categoryD1Ev _ZN12_GLOBAL__N_122generic_error_categoryD2Ev _ZN12_GLOBAL__N_122generic_error_categoryD1Ev _ZN12_GLOBAL__N_121system_error_categoryD0Ev _ZN12_GLOBAL__N_122generic_error_categoryD0Ev _ZNK12_GLOBAL__N_121system_error_category7messageEi _ZNK12_GLOBAL__N_122generic_error_category7messageEi _ZN12_GLOBAL__N_1L24system_category_instanceE _ZN12_GLOBAL__N_1L25generic_category_instanceE _GLOBAL__sub_I__ZNSt14error_categoryD2Ev _ZTSN12_GLOBAL__N_122generic_error_categoryE _ZTSN12_GLOBAL__N_121system_error_categoryE _ZTIN12_GLOBAL__N_121system_error_categoryE _ZTIN12_GLOBAL__N_122generic_error_categoryE _ZTVN12_GLOBAL__N_122generic_error_categoryE _ZTVN12_GLOBAL__N_121system_error_categoryE new_handler.cc _ZN12_GLOBAL__N_113__new_handlerE bad_array_new.cc cp-demangle.c d_make_comp d_make_name d_cv_qualifiers d_ref_qualifier d_substitution standard_subs d_count_templates_scopes d_append_char d_number.isra.0 d_number_component d_compact_number d_template_param d_discriminator d_source_name d_call_offset d_lookup_template_argument.isra.6 d_find_pack d_growable_string_callback_adapter d_append_string d_append_num d_print_comp d_print_expr_op d_print_subexpr cplus_demangle_builtin_types d_print_mod d_print_array_type.isra.10 d_print_function_type.isra.11 d_print_cast.isra.12 d_print_mod_list d_expr_primary d_type d_encoding d_template_args d_operator_name d_exprlist d_unqualified_name d_expression_1 d_vector_type d_function_type d_name d_parmlist d_bare_function_type cplus_demangle_operators d_demangle_callback.constprop.16 libgcc2.c unwind-dw2.c read_sleb128 execute_cfa_program uw_frame_state_for execute_stack_op dwarf_reg_size_table uw_update_context_1 uw_init_context_1 uw_update_context _Unwind_RaiseException_Phase2 _Unwind_ForcedUnwind_Phase2 uw_install_context_1 _Unwind_DebugHook .L18 .L97 .L208 .L294 .L485 .L20 .L21 .L22 .L23 .L24 .L25 .L26 .L27 .L28 .L29 .L30 .L31 .L32 .L33 .L34 .L35 .L36 .L37 .L38 .L39 .L40 .L41 .L42 .L43 .L61 .L55 .L56 .L62 .L59 .L60 .L183 .L177 .L178 .L184 .L181 .L182 .L217 .L211 .L212 .L218 .L215 .L216 .L303 .L297 .L298 .L299 .L300 .L301 .L305 .L306 .L307 .L308 .L309 .L310 .L311 .L312 .L313 .L314 .L315 .L316 .L317 .L318 .L319 .L320 .L321 .L402 .L323 .L341 .L335 .L336 .L342 .L339 .L340 .L378 .L380 .L381 .L382 .L383 .L384 .L385 .L386 .L387 .L388 .L389 .L390 .L391 .L392 .L393 .L394 .L395 .L486 .L488 .L489 .L490 .L491 unwind-dw2-fde.c fde_unencoded_compare frame_downheap frame_heapsort size_of_encoded_value base_from_object read_encoded_value_with_base fde_single_encoding_compare get_cie_encoding classify_object_over_fdes add_fdes linear_search_fdes fde_mixed_encoding_compare search_object terminator.6216 marker.6110 unseen_objects seen_objects .L80 .L89 .L83 .L84 .L90 .L87 .L88 /opt/MeetiXOSProject/MXlibraries/lib/crt0.o wait ps2_driver.cpp _ZStL19piecewise_construct _ZL20__gthread_key_deletei _ZStL8__ioinit _Z41__static_initialization_and_destruction_0ii _ZL16THREAD_TYPE_MAIN _ZL15THREAD_TYPE_SUB _ZL16THREAD_TYPE_VM86 _ZL22THREAD_PRIORITY_NORMAL _ZL20THREAD_PRIORITY_IDLE _ZL11FS_SEEK_SET _ZL11FS_SEEK_CUR _ZL11FS_SEEK_END _ZL17FS_NODE_TYPE_NONE _ZL17FS_NODE_TYPE_ROOT _ZL23FS_NODE_TYPE_MOUNTPOINT _ZL19FS_NODE_TYPE_FOLDER _ZL17FS_NODE_TYPE_FILE _ZL17FS_NODE_TYPE_PIPE _ZL34FS_REGISTER_AS_DELEGATE_SUCCESSFUL _ZL39FS_REGISTER_AS_DELEGATE_FAILED_EXISTING _ZL48FS_REGISTER_AS_DELEGATE_FAILED_DELEGATE_CREATION _ZL27FS_TRANSACTION_NO_REPEAT_ID _ZL22FS_TRANSACTION_WAITING _ZL23FS_TRANSACTION_FINISHED _ZL21FS_TRANSACTION_REPEAT _ZL29FS_CREATE_NODE_STATUS_CREATED _ZL29FS_CREATE_NODE_STATUS_UPDATED _ZL38FS_CREATE_NODE_STATUS_FAILED_NO_PARENT _ZL23FS_DISCOVERY_SUCCESSFUL _ZL22FS_DISCOVERY_NOT_FOUND _ZL17FS_DISCOVERY_BUSY _ZL18FS_DISCOVERY_ERROR _ZL40FS_TASKED_DELEGATE_REQUEST_TYPE_DISCOVER _ZL36FS_TASKED_DELEGATE_REQUEST_TYPE_READ _ZL37FS_TASKED_DELEGATE_REQUEST_TYPE_WRITE _ZL42FS_TASKED_DELEGATE_REQUEST_TYPE_GET_LENGTH _ZL46FS_TASKED_DELEGATE_REQUEST_TYPE_READ_DIRECTORY _ZL36FS_TASKED_DELEGATE_REQUEST_TYPE_OPEN _ZL37FS_TASKED_DELEGATE_REQUEST_TYPE_CLOSE _ZL18FS_OPEN_SUCCESSFUL _ZL17FS_OPEN_NOT_FOUND _ZL13FS_OPEN_ERROR _ZL12FS_OPEN_BUSY _ZL18FS_READ_SUCCESSFUL _ZL18FS_READ_INVALID_FD _ZL12FS_READ_BUSY _ZL13FS_READ_ERROR _ZL19FS_WRITE_SUCCESSFUL _ZL19FS_WRITE_INVALID_FD _ZL22FS_WRITE_NOT_SUPPORTED _ZL13FS_WRITE_BUSY _ZL14FS_WRITE_ERROR _ZL19FS_CLOSE_SUCCESSFUL _ZL19FS_CLOSE_INVALID_FD _ZL13FS_CLOSE_BUSY _ZL14FS_CLOSE_ERROR _ZL18FS_SEEK_SUCCESSFUL _ZL18FS_SEEK_INVALID_FD _ZL13FS_SEEK_ERROR _ZL18FS_TELL_SUCCESSFUL _ZL18FS_TELL_INVALID_FD _ZL20FS_LENGTH_SUCCESSFUL _ZL20FS_LENGTH_INVALID_FD _ZL19FS_LENGTH_NOT_FOUND _ZL14FS_LENGTH_BUSY _ZL15FS_LENGTH_ERROR _ZL21FS_CLONEFD_SUCCESSFUL _ZL28FS_CLONEFD_INVALID_SOURCE_FD _ZL16FS_CLONEFD_ERROR _ZL18FS_PIPE_SUCCESSFUL _ZL13FS_PIPE_ERROR _ZL32SET_WORKING_DIRECTORY_SUCCESSFUL _ZL34SET_WORKING_DIRECTORY_NOT_A_FOLDER _ZL31SET_WORKING_DIRECTORY_NOT_FOUND _ZL27SET_WORKING_DIRECTORY_ERROR _ZL32GET_WORKING_DIRECTORY_SUCCESSFUL _ZL35GET_WORKING_DIRECTORY_SIZE_EXCEEDED _ZL27GET_WORKING_DIRECTORY_ERROR _ZL28FS_OPEN_DIRECTORY_SUCCESSFUL _ZL27FS_OPEN_DIRECTORY_NOT_FOUND _ZL23FS_OPEN_DIRECTORY_ERROR _ZL28FS_READ_DIRECTORY_SUCCESSFUL _ZL21FS_READ_DIRECTORY_EOD _ZL23FS_READ_DIRECTORY_ERROR _ZL31FS_DIRECTORY_REFRESH_SUCCESSFUL _ZL26FS_DIRECTORY_REFRESH_ERROR _ZL25FS_DIRECTORY_REFRESH_BUSY _ZL26MESSAGE_SEND_MODE_BLOCKING _ZL30MESSAGE_SEND_MODE_NON_BLOCKING _ZL29MESSAGE_RECEIVE_MODE_BLOCKING _ZL33MESSAGE_RECEIVE_MODE_NON_BLOCKING _ZL30MESSAGE_SEND_STATUS_SUCCESSFUL _ZL30MESSAGE_SEND_STATUS_QUEUE_FULL _ZL26MESSAGE_SEND_STATUS_FAILED _ZL35MESSAGE_SEND_STATUS_EXCEEDS_MAXIMUM _ZL33MESSAGE_RECEIVE_STATUS_SUCCESSFUL _ZL34MESSAGE_RECEIVE_STATUS_QUEUE_EMPTY _ZL29MESSAGE_RECEIVE_STATUS_FAILED _ZL43MESSAGE_RECEIVE_STATUS_FAILED_NOT_PERMITTED _ZL42MESSAGE_RECEIVE_STATUS_EXCEEDS_BUFFER_SIZE _ZL34MESSAGE_RECEIVE_STATUS_INTERRUPTED _ZL26EVAQUERY_STATUS_SUCCESSFUL _ZL26EVAQUERY_STATUS_UNKNOWN_ID _GLOBAL__sub_I_mousePacketNumber ps2_driver_irq_triggered.cpp _GLOBAL__sub_I__Z21registerOperationModev ps2_driver_polling.cpp _GLOBAL__sub_I_ps2_driver_polling.cpp flog.cpp _GLOBAL__sub_I__ZN7FileLog4flogESs logger.cpp utils.cpp eh_term_handler.cc eh_unex_handler.cc globals_io.cc AllocMem.cpp AtomicBlock.cpp GetPidForTid.cpp GetTid.cpp GetWorkingDirectory.cpp Log.cpp ReceiveMessage.cpp RegisterIrqHandler.cpp RestoreInterruptedState.cpp SendMessage.cpp SetWorkingDirectory.cpp ShareMem.cpp syscall.cpp TaskRegisterID.cpp __AtomicLock.cpp isalnum.cpp isalpha.cpp iscntrl.cpp isgraph.cpp islower.cpp isprint.cpp ispunct.cpp isspace.cpp isupper.cpp isxdigit.cpp tolower.cpp toupper.cpp errno.cpp itanium_cxx_abi_support.cpp setlocale.cpp main.cpp dlmalloc.cpp _ZL17spin_acquire_lockPi _ZL19malloc_global_mutex _ZL7mparams _ZL4_gm_ _ZL15segment_holdingP12malloc_statePc _ZL16has_segment_linkP12malloc_stateP14malloc_segment _ZL12init_mparamsv _ZL13change_mparamii _ZL17internal_mallinfoP12malloc_state _ZL21internal_malloc_statsP12malloc_state _ZL10mmap_allocP12malloc_statem _ZL11mmap_resizeP12malloc_stateP12malloc_chunkmi _ZL8init_topP12malloc_stateP12malloc_chunkm _ZL9init_binsP12malloc_state _ZL13prepend_allocP12malloc_statePcS1_m _ZL11add_segmentP12malloc_statePcmj _ZL9sys_allocP12malloc_statem _ZL23release_unused_segmentsP12malloc_state _ZL8sys_trimP12malloc_statem _ZL13dispose_chunkP12malloc_stateP12malloc_chunkm _ZL13tmalloc_largeP12malloc_statem _ZL13tmalloc_smallP12malloc_statem _ZL17try_realloc_chunkP12malloc_stateP12malloc_chunkmi _ZL17internal_memalignP12malloc_statemm _ZL6iallocP12malloc_statemPmiPPv _ZL18internal_bulk_freeP12malloc_statePPvm sched_yield.cpp signal.cpp fclose.cpp __fclose_static.cpp __fclose_static_unlocked.cpp fdopen.cpp __fdopen_static.cpp fflush.cpp __fflush_unlocked.cpp __fflush_write_unlocked.cpp fileno.cpp fopen.cpp __fopen_static.cpp fprintf.cpp fputc.cpp __fputc_unlocked.cpp fputs.cpp fread.cpp __fread_unlocked.cpp fseek.cpp __fseeko_unlocked.cpp ftell.cpp __ftello_unlocked.cpp fwrite.cpp __fwrite_unlocked.cpp getc.cpp __open_file_list.cpp __parse_mode_flags.cpp putc.cpp __setdefbuf_unlocked.cpp setvbuf.cpp __setvbuf_unlocked.cpp sprintf.cpp sscanf.cpp stdio.cpp __stdio_impl_close.cpp __stdio_impl_eof.cpp __stdio_impl_error.cpp __stdio_impl_fileno.cpp __stdio_impl_read.cpp __stdio_impl_reopen.cpp __stdio_impl_seek.cpp __stdio_impl_tell.cpp __stdio_impl_write.cpp ungetc.cpp vfprintf.cpp __vfprintf_unlocked.cpp _ZL27vcbprintf_vfprintf_callbackPvPKcm vsnprintf.cpp _ZL28vcbprintf_vsnprintf_callbackPvPKcm vsprintf.cpp abort.cpp exit.cpp parseargs.cpp strtod.cpp strtof.cpp memchr.cpp memcmp.cpp memcpy.cpp memmove.cpp memset.cpp strcmp.cpp strcoll.cpp strcpy.cpp strerror.cpp strlen.cpp strxfrm.cpp fstat.cpp strftime.cpp time.cpp close.cpp lseek.cpp read.cpp sbrk.cpp tell.cpp write.cpp open.cpp basename.cpp _ZL8_statbuf sig_handlers.cpp __fflush_read_unlocked.cpp __fgetc_unlocked.cpp __fungetc_unlocked.cpp klog.cpp kvlog.cpp vcbprintf.cpp _ZL11_get_numberPPKc _ZL18_integer_to_stringPcyyPKc strncpy.cpp strrchr.cpp AtomicLock.cpp AtomicTryLock.cpp CliArgsRelease.cpp Close.cpp Exit.cpp GetExecutablePath.cpp Millis.cpp Open.cpp Read.cpp RegisterSignalHandler.cpp Sbrk.cpp Seek.cpp Tell.cpp Write.cpp Yield.cpp _GLOBAL_OFFSET_TABLE_ __x86.get_pc_thunk.cx _ZNSo5writeEPKcl _ZNSs2atEm _ZNSt10ctype_base5digitE __cxa_free_exception _ZNSirsERf _ZNSsC1IN9__gnu_cxx17__normal_iteratorIPcSsEEEET_S4_RKSaIcE _ZNSt13basic_fstreamIcSt11char_traitsIcEE7is_openEv _ZNSirsERj _ZTSSt18basic_stringstreamIcSt11char_traitsIcESaIcEE _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_PS3_ _ZNKSt9type_info15__is_function_pEv _ZTVN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE _ZSt10unexpectedv _ZNSt6localeC2EPNS_5_ImplE _ZTTSt14basic_ifstreamIcSt11char_traitsIcEE _ZNSolsEPSt15basic_streambufIcSt11char_traitsIcEE _ZSt18__throw_bad_typeidv _ZNKSt11__timepunctIcE7_M_daysEPPKc _ZNSaIwEC1Ev _ZNSt14overflow_errorC1ERKSs _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb _ZTSSt19basic_ostringstreamIcSt11char_traitsIcESaIcEE strcpy _ZNSt9basic_iosIcSt11char_traitsIcEEC2Ev _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm Tell _ZNKSs6substrEmm _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecm __main _ZNSt17moneypunct_bynameIcLb0EE4intlE _ZTCSd0_Si _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Em _stdin_buf _Unwind_Find_FDE realloc_in_place _ZN10__cxxabiv115__forced_unwindD1Ev _ZNSt14codecvt_bynameIcc9mbstate_tED2Ev _ZNSs4nposE _ZNKSt5ctypeIcE8do_widenEPKcS2_Pc _ZNSt15basic_streambufIcSt11char_traitsIcEE5sputnEPKcl _ZNSt8messagesIcE2idE _ZNSt16__numpunct_cacheIcED2Ev _ZNSt9basic_iosIcSt11char_traitsIcEE4initEPSt15basic_streambufIcS1_E _Unwind_GetIPInfo _ZTSNSt6locale5facetE _ZNSt12__basic_fileIcE7seekoffExSt12_Ios_Seekdir _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKc _ZTVSt15messages_bynameIcE _ZNSt6locale13_S_initializeEv __cxa_demangle _ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Rh _ZTVSd _ZNSi10_M_extractImEERSiRT_ _ZNKSt13basic_fstreamIcSt11char_traitsIcEE7is_openEv _ZNSt17moneypunct_bynameIcLb1EEC2EPKcm _ZTVSt17bad_function_call __cxa_rethrow _ZNKSt15basic_streambufIcSt11char_traitsIcEE5ebackEv _ZTISt21__ctype_abstract_baseIcE _ZNKSs6rbeginEv _ZNSt10moneypunctIcLb0EED2Ev _ZSt14set_unexpectedPFvvE _ZNKSt10moneypunctIcLb0EE13do_neg_formatEv mousePacketNumber _ZTv0_n12_NSt13basic_fstreamIcSt11char_traitsIcEED1Ev _ZNSi5seekgESt4fposI9mbstate_tE _ZNSs12_S_constructIN9__gnu_cxx17__normal_iteratorIPcSsEEEES2_T_S4_RKSaIcESt20forward_iterator_tag __AtomicLock _ZNSs13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIS_SsEES2_ _ZTv0_n12_NSt14basic_ofstreamIcSt11char_traitsIcEED0Ev _ZNSs7replaceEmmRKSs _Unwind_GetIP _ZNSt6locale5facet17_S_clone_c_localeERPi _ZNSt14basic_ofstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode _ZNSoD1Ev _ZNSt12length_errorC1ERKSs _ZNSolsEl _ZNKSt5ctypeIcE5widenEPKcS2_Pc _ZNSt13basic_fstreamIcSt11char_traitsIcEEC1Ev _ZNSt15basic_streambufIcSt11char_traitsIcEED0Ev _ZNSs5beginEv _ZNSt9bad_allocD2Ev _ZNSt15basic_streambufIcSt11char_traitsIcEED1Ev stdout _ZNKSs5crendEv _ZTTSt19basic_istringstreamIcSt11char_traitsIcESaIcEE vsprintf _ZNSi5ungetEv _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEESt16initializer_listIcE _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEED0Ev _ZNK10__cxxabiv120__si_class_type_info20__do_find_public_srcElPKvPKNS_17__class_type_infoES2_ _ZNSt15basic_streambufIcSt11char_traitsIcEE9pbackfailEi _ZNSt6locale10_S_classicE _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_bRSt8ios_basecRKSs Yield _ZNSt10moneypunctIcLb0EE24_M_initialize_moneypunctEPiPKc _ZNSt6localeC1ERKS_ _ZTSSt14overflow_error _ZNKSs4backEv _ZTVNSt6locale5facetE _ZNSt5ctypeIcEC2EPKjbm _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecPKv _ZNSolsEy _ZNSt14collate_bynameIcED1Ev _ZTISt15basic_streambufIcSt11char_traitsIcEE __cxa_free_dependent_exception _ZNSt6locale5facetD0Ev _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED0Ev _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEEC2ESt13_Ios_Openmode _ZNSt12__basic_fileIcEC1EPi _ZNSs6assignEPKcm _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm __register_frame _ZN10__cxxabiv120__si_class_type_infoD2Ev _ZTSN10__cxxabiv120__si_class_type_infoE _ZTVSo _ZTSSt10moneypunctIcLb1EE _ZSt9has_facetISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZNSt8ios_base6badbitE ungetc _ZNKSt11__timepunctIcE19_M_days_abbreviatedEPPKc vcbprintf _ZNSt6locale5facet13_S_get_c_nameEv _ZNSt13basic_filebufIcSt11char_traitsIcEE27_M_allocate_internal_bufferEv _ZNSt12future_errorD1Ev _ZNKSt7collateIcE7compareEPKcS2_S2_S2_ _ZNSs7_M_moveEPcPKcm _ZN10__cxxabiv115__forced_unwindD2Ev _ZNK10__cxxabiv121__vmi_class_type_info11__do_upcastEPKNS_17__class_type_infoEPKvRNS1_15__upcast_resultE _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt8ios_base9showpointE _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Em _ZSt20__throw_future_errori _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv _ZSt2wsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_ _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKc _ZNSt9basic_iosIcSt11char_traitsIcEEC1EPSt15basic_streambufIcS1_E _ZSt18uncaught_exceptionv _ZSt9use_facetISt10moneypunctIcLb0EEERKT_RKSt6locale __open_file_list_remove _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St5_Setw _ZTISt15underflow_error _ZSt16__convert_from_vRKPiPciPKcz strerror _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEEC2ESt13_Ios_Openmode _ZTISt23__codecvt_abstract_baseIcc9mbstate_tE _ZNSt11__timepunctIcED2Ev _ZNSsD2Ev _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St14_Resetiosflags _ZNSt16__numpunct_cacheIcED0Ev __cxa_deleted_virtual _ZTCSt19basic_ostringstreamIcSt11char_traitsIcESaIcEE0_So _ZNSt13basic_filebufIcSt11char_traitsIcEEC1Ev _ZNSspLEc _ZNSt14basic_ofstreamIcSt11char_traitsIcEE7is_openEv _ZNSs6appendEmc _ZNSiD0Ev _ZSt19__throw_regex_errorNSt15regex_constants10error_typeE _ZNSt15basic_streambufIcSt11char_traitsIcEE6sbumpcEv memmove _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED2Ev _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_RS3_ _ZTVSt17moneypunct_bynameIcLb0EE _ZNSt17moneypunct_bynameIcLb1EED1Ev _ZNSt10moneypunctIcLb0EEC1EPiPKcm _ZNKSt15basic_streambufIcSt11char_traitsIcEE5egptrEv _ZTVSt10moneypunctIcLb1EE _ZNSt9exceptionD2Ev _Unwind_Resume_or_Rethrow syscall _ZTTSo _ZTVSt13basic_filebufIcSt11char_traitsIcEE _ZNSolsEb _ZNSs13_S_copy_charsEPcN9__gnu_cxx17__normal_iteratorIPKcSsEES4_ _ZNSt10ctype_base5spaceE _ZTISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZNKSt14basic_ofstreamIcSt11char_traitsIcEE7is_openEv _ZNKSt10moneypunctIcLb1EE11curr_symbolEv _ZTSSt12out_of_range _ZNSt8ios_base10floatfieldE _ZTISt8bad_cast _ZNSo9_M_insertIxEERSoT_ __fopen_static _ZNSs7_M_copyEPcPKcm _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl _ZNSsaSEPKc _Z12writeToMouseh _ZGVNSt8messagesIcE2idE _ZNSt15messages_bynameIcED2Ev AtomicTryLock GetWorkingDirectoryL _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC2EP4FILE _ZSt19__throw_ios_failurePKc _ZTISt8ios_base _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_bRSt8ios_basece _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZTVSt13bad_exception _ZSt17__copy_streambufsIcSt11char_traitsIcEElPSt15basic_streambufIT_T0_ES6_ _ZNSt20bad_array_new_lengthD1Ev _ZNSt12system_errorD2Ev _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt14overflow_errorD0Ev _ZTVSt8messagesIcE _ZTVSt11regex_error ReceiveMessage GetWorkingDirectory malloc_stats _ZNKSt15basic_streambufIcSt11char_traitsIcEE5pbaseEv _ZNSt6locale3allE _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE9underflowEv _ZNSt6locale5facetD1Ev _ZTVSt19basic_ostringstreamIcSt11char_traitsIcESaIcEE _ZTISt10ctype_base _ZNSs4_Rep11_S_terminalE _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt6locale5_Impl16_M_replace_facetEPKS0_PKNS_2idE _ZTSSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZGVNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZN5Utils12outportShortEtt _ZNKSs16find_last_not_ofEPKcmm _ZNSt14codecvt_bynameIcc9mbstate_tED1Ev _ZNSt14overflow_errorD2Ev _ZTISt18__moneypunct_cacheIcLb1EE __fungetc_unlocked _ZNSt18__moneypunct_cacheIcLb0EEC1Em _Unwind_GetRegionStart _ZNSt10ctype_base5graphE _ZNSt8ios_base7showposE _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intImEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNSt6locale5facet20_S_lc_ctype_c_localeEPiPKc irqHandler Write _ZNSt17moneypunct_bynameIcLb0EEC1EPKcm _ZNSt13basic_filebufIcSt11char_traitsIcEE9showmanycEv _ZNSt13basic_filebufIcSt11char_traitsIcEE5closeEv _ZNSt12out_of_rangeD2Ev _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev Read _ZNSt10moneypunctIcLb1EE4intlE _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED2Ev _ZTSSt19basic_istringstreamIcSt11char_traitsIcESaIcEE _ZNSdC1Ev _Znwm _ZNSt12system_errorD1Ev _ZNSt12future_errorD0Ev _ZNSs4_Rep10_M_disposeERKSaIcE __setvbuf_unlocked errno _ZNSiC2EPSt15basic_streambufIcSt11char_traitsIcEE __cxa_throw_bad_array_length _ZNKSt7collateIcE10_M_compareEPKcS2_ _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSs _ZNSsC2EmcRKSaIcE _ZNSt6locale5_ImplD1Ev _ZNSt15basic_streambufIcSt11char_traitsIcEE9showmanycEv keyboardReceiverTid _ZNSt6locale5_Impl11_S_id_ctypeE _ZNSsC1ERKSs _ZNKSs7compareEPKc _ZNKSt9basic_iosIcSt11char_traitsIcEE6narrowEcc _ZNSt11__timepunctIcEC2Em _ZNKSt19basic_ostringstreamIcSt11char_traitsIcESaIcEE3strEv _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRSs _ZTv0_n12_NSt14basic_ofstreamIcSt11char_traitsIcEED1Ev _ZNSt15basic_streambufIcSt11char_traitsIcEE12__safe_gbumpEl _ZSt13__int_to_charIcyEiPT_T0_PKS0_St13_Ios_Fmtflagsb _Unwind_Backtrace _ZNKSt5ctypeIcE10do_tolowerEPcPKc _ZNKSt7codecvtIcc9mbstate_tE16do_always_noconvEv _ZNKSs4copyEPcmm _ZNSt8ios_base6eofbitE _ZTVSt18__moneypunct_cacheIcLb1EE _ZNSt11regex_errorD1Ev _ZNSt6localeC1Ev Open _ZNKSt10error_code23default_error_conditionEv _ZNSt8ios_base3outE Sbrk _ZNSirsERm _ZNSt16__numpunct_cacheIcED1Ev _ZNKSt10moneypunctIcLb1EE13do_pos_formatEv _ZNSt10bad_typeidD0Ev _ZNSt15basic_streambufIcSt11char_traitsIcEEC1ERKS2_ _ZNSt14overflow_errorD1Ev _ZNSo5flushEv _ZNSt8messagesIcED1Ev _ZNSt7collateIcED0Ev _ZNKSt10moneypunctIcLb0EE16do_decimal_pointEv _ZNSt12__basic_fileIcE8xsputn_2EPKclS2_l _ZNKSt8numpunctIcE8groupingEv _ZNKSt10moneypunctIcLb0EE10neg_formatEv _ZNSt8bad_castD0Ev _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy _ZNSaIwED1Ev _ZNSt8ios_baseD1Ev _ZNSs6assignEmc _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNSt15basic_streambufIcSt11char_traitsIcEE5sgetnEPcl _ZNKSs4_Rep12_M_is_leakedEv _ZTVSt13basic_fstreamIcSt11char_traitsIcEE _ZNSt10ctype_base6xdigitE _stderr __cxa_call_unexpected _ZNSt15basic_streambufIcSt11char_traitsIcEEC1Ev _ZNKSt10moneypunctIcLb1EE16do_positive_signEv _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4fileEv _ZNSt13basic_filebufIcSt11char_traitsIcEE5imbueERKSt6locale _ZNSi10_M_extractItEERSiRT_ __cxa_get_exception_ptr _ZNSi10_M_extractIdEERSiRT_ _ZTISd _ZSt4cerr _ZNSdD1Ev _ZNSt10moneypunctIcLb0EEC2Em _ZNSsC2ESt16initializer_listIcERKSaIcE _ZNSt12__basic_fileIcE2fdEv _ZNSt6locale5_ImplC1Em _ZNKSsixEm _ZNKSt13basic_filebufIcSt11char_traitsIcEE7is_openEv _ZNSt12length_errorD2Ev _ZNSolsEt _ZN6Logger3logEPKcz _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRb _ZNSt8ios_base17register_callbackEPFvNS_5eventERS_iEi _ZSt9has_facetISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZNKSt10moneypunctIcLb1EE10pos_formatEv RestoreInterruptedState _ZNSirsERi _ZNKSt7collateIcE10do_compareEPKcS2_S2_S2_ _ZNSirsEPFRSt9basic_iosIcSt11char_traitsIcEES3_E _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intImEES3_S3_RSt8ios_basecT_ _ZTISt15basic_stringbufIcSt11char_traitsIcESaIcEE _ZNSt10moneypunctIcLb1EEC1EPiPKcm _ZNSt13basic_fstreamIcSt11char_traitsIcEEC2Ev _ZNSt15messages_bynameIcEC2EPKcm getc _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecx _ZTVSt12out_of_range _ZNSt6locale5_ImplC2Em _Unwind_GetCFA _ZSt13set_terminatePFvvE memcpy _ZNKSt15basic_stringbufIcSt11char_traitsIcESaIcEE3strEv _ZNSsC2Ev _ZTSSt14basic_ifstreamIcSt11char_traitsIcEE _ZNSt14basic_ifstreamIcSt11char_traitsIcEE7is_openEv _ZNSt17__timepunct_cacheIcEC2Em _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Em _ZNKSs17find_first_not_ofERKSsm _ZNKSs17find_first_not_ofEPKcmm _ZNKSt7collateIcE12do_transformEPKcS2_ setvbuf __cxa_allocate_dependent_exception __TMC_END__ _ZTISt15numpunct_bynameIcE _ZTVSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZNSt6locale5facet19_S_destroy_c_localeERPi _ZNSsC1IPKcEET_S2_RKSaIcE _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_c _ZTVSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZTVSt23__codecvt_abstract_baseIcc9mbstate_tE _ZSt9has_facetISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale open_file_list_lockatom SendMessage _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basece _ZNKSt10moneypunctIcLb1EE16do_thousands_sepEv _ZTVSt11range_error _ZNKSt8messagesIcE4openERKSsRKSt6localePKc _ZNSt13runtime_errorD2Ev _ZNSt7codecvtIcc9mbstate_tEC1EPim _ZTCSt14basic_ofstreamIcSt11char_traitsIcEE0_So _ZNSt10moneypunctIcLb0EE2idE _ZSt21__throw_runtime_errorPKc __stdio_impl_error _ZNSt17__timepunct_cacheIcE12_S_timezonesE __DTOR_END__ _ZNSt13basic_fstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode _ZNKSs5rfindEPKcm _ZN9__gnu_cxx4ropeIcSaIcEE10_S_min_lenE _ZTISt10money_base _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6_M_padEclRSt8ios_basePcPKcRi _ZTVSt16invalid_argument _ZN10__cxxabiv117__class_type_infoD1Ev _ZNSt11logic_errorC2ERKSs _ZTVSt14basic_ifstreamIcSt11char_traitsIcEE _ZN9__gnu_cxxeqIPKcSsEEbRKNS_17__normal_iteratorIT_T0_EES8_ _ZTIN10__cxxabiv121__vmi_class_type_infoE _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_EPKS3_RKS6_ _ZNSt13basic_filebufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZNSaIcED2Ev _ZNSirsERd _ZTSSt12codecvt_base _ZTVSt11__timepunctIcE _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE7seekposESt4fposI9mbstate_tESt13_Ios_Openmode islower _ZNKSt11__timepunctIcE15_M_time_formatsEPPKc _ZNSt7codecvtIcc9mbstate_tEC2EPim _ZTSSt17moneypunct_bynameIcLb0EE _ZNSt11range_errorC2ERKSs _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEE3strERKSs _ZNSi7putbackEc tolower _ZNSt13basic_filebufIcSt11char_traitsIcEE15_M_create_pbackEv _ZNSt15messages_bynameIcEC1EPKcm _ZNSt7collateIcEC1EPim _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcm _ZNSsaSERKSs _ZTIN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEE _ZNSt6locale18_S_initialize_onceEv _ZTISt12out_of_range _ZNKSs15_M_check_lengthEmmPKc _ZNSt10ctype_base5printE _ZTSSt14collate_bynameIcE _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Em _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNSs12_S_constructEmcRKSaIcE _ZNSt10__num_base15_S_format_floatERKSt8ios_basePcc _ZNSaIcEC1Ev _ZNSt20bad_array_new_lengthD2Ev _ZNKSt7codecvtIcc9mbstate_tE6do_outERS0_PKcS4_RS4_PcS6_RS6_ malloc _ZTSSt20bad_array_new_length _ZNKSt11__timepunctIcE8_M_am_pmEPPKc _ZNSt8messagesIcEC1Em _ZNSi6sentryC2ERSib _ZNSi3getEPclc _ZNSt15basic_streambufIcSt11char_traitsIcEE5gbumpEi _ZTSSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZNSo3putEc _ZTVSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZNSs15_M_replace_safeEmmPKcm _ZSt22__throw_overflow_errorPKc _ZNSolsEf OpenF _ZNSt13basic_filebufIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode _ZTVSt7codecvtIcc9mbstate_tE _ZNKSt6localeeqERKS_ OpenFMS _ZNSt9basic_iosIcSt11char_traitsIcEE7copyfmtERKS2_ _ZNSt6locale5_Impl16_M_install_facetEPKNS_2idEPKNS_5facetE _ZNSt18__moneypunct_cacheIcLb1EED0Ev _ZNSt12out_of_rangeC2ERKSs _ZNSt7collateIcED2Ev _ZNSt6locale5_ImplD2Ev _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_h _ZNSo6sentryD2Ev vsnprintf _ZTSSt16__numpunct_cacheIcE _ZNSi10_M_extractIeEERSiRT_ _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1ERKSsSt13_Ios_Openmode _ZNSt15basic_streambufIcSt11char_traitsIcEE5pbumpEi _ZNSs7reserveEm _ZNKSs7compareEmmPKc _ZTTSt19basic_ostringstreamIcSt11char_traitsIcESaIcEE SeekS _ZSt15system_categoryv _ZGVNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNKSs4sizeEv _ZNSs9_M_mutateEmmm _ZNSs7replaceEmmPKcm _ZNKSs16find_last_not_ofEcm _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE3strERKSs _ZNSt15numpunct_bynameIcED0Ev _ZNSolsEm _ZNSt7codecvtIcc9mbstate_tED0Ev _ZNSt6locale5_Impl13_S_id_numericE _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKcm _ZNSt6locale5_ImplC2ERKS0_m _ZNKSt5ctypeIcE13_M_widen_initEv __dso_handle _ZNSs6appendEPKc _ZNSt14basic_ifstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode _ZNSt10__num_base11_S_atoms_inE _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode _ZTSSt8ios_base SendMessageT _ZNKSt10moneypunctIcLb0EE10pos_formatEv _ZN10__cxxabiv121__vmi_class_type_infoD1Ev __stdio_impl_reopen _ZNKSs17find_first_not_ofEcm _ZNK10__cxxabiv117__class_type_info10__do_catchEPKSt9type_infoPPvj _ZNSi6ignoreEv _ZNSt8ios_base4InitC2Ev _ZNKSs9_M_ibeginEv _ZNSt12__basic_fileIcE4fileEv _ZNSt13runtime_errorC2ERKSs _ZNKSt10moneypunctIcLb0EE14do_curr_symbolEv _ZNSt9basic_iosIcSt11char_traitsIcEE11_M_setstateESt12_Ios_Iostate _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecb ispunct _ZTCSt13basic_fstreamIcSt11char_traitsIcEE0_Sd _ZNSt10moneypunctIcLb1EEC2Em _ZNSt13basic_filebufIcSt11char_traitsIcEE4openERKSsSt13_Ios_Openmode __stdio_impl_read _ZNSt8ios_base6skipwsE _ZNSt17moneypunct_bynameIcLb0EED2Ev _ZNSi3getEPcl _ZNKSt10moneypunctIcLb1EE11frac_digitsEv _ZN7FileLog4flogESs _ZNSt8numpunctIcED0Ev _ZTSSo _ZNSt12__basic_fileIcE4openEPKcSt13_Ios_Openmodei _ZTVSt9type_info _ZTTSt14basic_ofstreamIcSt11char_traitsIcEE _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZTSSt16invalid_argument _ZNSt6locale5_Impl19_S_facet_categoriesE _ZSt17__throw_bad_allocv _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2Ev _ZZNSt13basic_filebufIcSt11char_traitsIcEE5closeEvEN14__close_sentryD2Ev _ZNSt13basic_filebufIcSt11char_traitsIcEE14_M_get_ext_posER9mbstate_t __frame_state_for SetWorkingDirectory _ZNSt15basic_streambufIcSt11char_traitsIcEE8overflowEi _ZNSt13basic_fstreamIcSt11char_traitsIcEE4openEPKcSt13_Ios_Openmode _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC2Em _ZTSSt8messagesIcE malloc_footprint_limit _ZNSirsERt _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Em _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNKSt9exception4whatEv _ZNKSs4findEcm _ZNSaIwEC2Ev pvalloc _ZNKSs16find_last_not_ofEPKcm _ZTVSt16bad_array_length _ZTSSt18__moneypunct_cacheIcLb0EE isspace _ZNSt8numpunctIcEC2EPSt16__numpunct_cacheIcEm _ZNKSs4findEPKcm _stdin _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt _ZNKSs12find_last_ofEPKcm _ZTISt11regex_error _ZTSSt13basic_filebufIcSt11char_traitsIcEE _ZNKSs5rfindEPKcmm _ZNKSt8messagesIcE8do_closeEi _ZTISt9bad_alloc _ZNSt13basic_filebufIcSt11char_traitsIcEE4syncEv _ZNKSs6_M_repEv fflush _ZSt16generic_categoryv _ZTSSt7collateIcE _ZNSt6locale5_Impl14_S_id_monetaryE _ZTCSt18basic_stringstreamIcSt11char_traitsIcESaIcEE8_So _ZNKSt19basic_ostringstreamIcSt11char_traitsIcESaIcEE5rdbufEv __fread_unlocked _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE8overflowEi _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf _ZNSs5eraseEN9__gnu_cxx17__normal_iteratorIPcSsEE _ZN14__gnu_internal8buf_cerrE _ZSt9use_facetISt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZNSt6locale4timeE _ZNSt13basic_filebufIcSt11char_traitsIcEE19_M_terminate_outputEv _ZSt9use_facetISt8numpunctIcEERKT_RKSt6locale _ZNKSt10moneypunctIcLb1EE13thousands_sepEv _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE21_M_extract_via_formatES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tmPKc _ZSt9has_facetISt7codecvtIcc9mbstate_tEEbRKSt6locale _ZNSs6assignERKSs _ZN5Utils11inportShortEt _ZNSsixEm _ZGVNSt11__timepunctIcE2idE _ZTVSt18basic_stringstreamIcSt11char_traitsIcESaIcEE TaskRegisterID _FiniLibc _ZNSt8numpunctIcEC1Em _ZTVSt8ios_base _ZTISt17bad_function_call _ZNSs6assignEOSs _ZN14__gnu_internal13buf_cerr_syncE _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_bRSt8ios_basece _ZSt14__convert_to_vIfEvPKcRT_RSt12_Ios_IostateRKPi _ZTSSt8numpunctIcE _ZTVN10__cxxabiv120__si_class_type_infoE _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St8_Setbase _ZGVNSt7collateIcE2idE _ZSt9use_facetISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZThn8_NSdD0Ev _ZNSsD1Ev _ZNSolsEPFRSoS_E _ZNSt8bad_castD1Ev __umoddi3 lseek _ZTSSt10money_base _ZNSs3endEv independent_calloc _ZNSt9basic_iosIcSt11char_traitsIcEED2Ev _ZTVSt11logic_error _ZNK10__cxxabiv117__class_type_info11__do_upcastEPKS0_PKvRNS0_15__upcast_resultE _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE9pbackfailEi _ZdlPv _ZNSt13basic_filebufIcSt11char_traitsIcEE6xsputnEPKcl _ZN9__gnu_cxx20recursive_init_errorD1Ev _ZNSi4peekEv _ZNSt8messagesIcEC2Em _ZNSt12length_errorD0Ev _ZSt9use_facetISt11__timepunctIcEERKT_RKSt6locale _ZNSt10money_base18_S_default_patternE _ZN10__cxxabiv121__vmi_class_type_infoD0Ev _ZNSt10ctype_base5lowerE _ZNSt8ios_base6binaryE _ZSt15get_new_handlerv _ZTISt15messages_bynameIcE _ZNSt18__moneypunct_cacheIcLb1EEC2Em _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEED1Ev _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEEC2ESt13_Ios_Openmode _ZNSo6sentryD1Ev __udivdi3 _ZNSt15basic_streambufIcSt11char_traitsIcEE6xsputnEPKcl _ZTVSt14overflow_error _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcm _ZNSt8ios_base5imbueERKSt6locale _ZSt20__throw_length_errorPKc __fgetc_unlocked _ZTSSt14error_category _ZNSi7getlineEPcl abort _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1Ev _ZNSt15basic_streambufIcSt11char_traitsIcEE9pubsetbufEPcl _ZNSolsEPKv _ZNSt17moneypunct_bynameIcLb1EE4intlE _ZSt14__add_groupingIcEPT_S1_S0_PKcmPKS0_S5_ _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE4syncEv _ZNKSt9basic_iosIcSt11char_traitsIcEE3eofEv _ZNSs4_Rep10_M_refcopyEv _ZTVSi _ZNKSt11__use_cacheISt16__numpunct_cacheIcEEclERKSt6locale _ZSt17__verify_groupingPKcmRKSs _ZNSirsEPSt15basic_streambufIcSt11char_traitsIcEE _ZNSt15basic_streambufIcSt11char_traitsIcEE6setbufEPcl _ZNSt10ctype_base5alphaE _ZNSs18_S_construct_aux_2EmcRKSaIcE GetPidForTid _ZTCSt13basic_fstreamIcSt11char_traitsIcEE0_Si sig_handler_SIG_IGN __cxa_end_catch _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEEC2ERKSsSt13_Ios_Openmode _ZTISt9basic_iosIcSt11char_traitsIcEE isxdigit _ZNSt12__basic_fileIcE6xsgetnEPcl _ZTISo _ZNKSt7codecvtIcc9mbstate_tE10do_unshiftERS0_PcS3_RS3_ _ZNSt13bad_exceptionD2Ev _init _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZN5Utils9inportIntEt _ZNSsC1ESt16initializer_listIcERKSaIcE _ZTSSt12system_error _ZN14__gnu_internal7buf_cinE ReceiveMessageTMB _ZNSt14codecvt_bynameIcc9mbstate_tEC2EPKcm _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt8ios_base3begE _ZNKSt7collateIcE9transformEPKcS2_ _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St8_Setbase _ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Pa _ZNSt15basic_streambufIcSt11char_traitsIcEE6xsgetnEPcl _ZNKSs4_Rep12_M_is_sharedEv _ZNSt9basic_iosIcSt11char_traitsIcEE5imbueERKSt6locale _ZNKSt5ctypeIcE10do_toupperEPcPKc _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKh _ZNKSt10moneypunctIcLb0EE13positive_signEv _ZNKSs7_M_dataEv _ZNSt17moneypunct_bynameIcLb1EED0Ev _ZNSsC2ERKSsmmRKSaIcE _ZNKSt6locale4nameEv _ZNSt12__basic_fileIcED1Ev _ZSt9terminatev _ZNSs6resizeEm _ZNSi6ignoreEli _ZNSo9_M_insertIeEERSoT_ _ZNSaIcEC2ERKS_ _ZSt24__throw_out_of_range_fmtPKcz _ZNSt15underflow_errorD1Ev _ZNSt10money_base20_S_construct_patternEccc _ZTSSt12future_error _ZNSt13basic_fstreamIcSt11char_traitsIcEED0Ev _ZSt24__throw_invalid_argumentPKc _ZNSs6assignEPKc _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRf _ZNSs4_Rep7_M_grabERKSaIcES2_ _ZNSs6insertEmRKSsmm _ZNKSt10moneypunctIcLb0EE13decimal_pointEv _ZNSt6locale5facet18_S_initialize_onceEv bulk_free _ZNKSs5frontEv __register_frame_table _ZNKSt8ios_base7failure4whatEv _ZNSt8ios_base20_M_dispose_callbacksEv _ZNSt11logic_errorD0Ev _ZNSt17moneypunct_bynameIcLb1EED2Ev _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEEC1ESt13_Ios_Openmode _ZN10__cxxabiv119__foreign_exceptionD2Ev _ZNSt14collate_bynameIcEC2EPKcm _ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPK2tmPKcSB_ _ZNKSs13find_first_ofEPKcm _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2Em _ZNKSt5ctypeIcE10do_tolowerEc _ZNSt5ctypeIcEC1EPiPKjbm _ZSt7getlineIcSt11char_traitsIcESaIcEERSt13basic_istreamIT_T0_ES7_RSbIS4_S5_T1_ES4_ _ZNSt6locale5_Impl16_M_install_cacheEPKNS_5facetEm _ZTSN10__cxxabiv117__class_type_infoE _ZTSSt23__codecvt_abstract_baseIcc9mbstate_tE strrchr _ZSt9has_facetISt10moneypunctIcLb0EEEbRKSt6locale _ZNSirsEPFRSiS_E _ZNSt8ios_base7failbitE basename _ZTISt9time_base _ZNSs6appendERKSsmm _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE14_M_group_floatEPKcmcS6_PcS7_Ri _ZNSt18__moneypunct_cacheIcLb0EE8_M_cacheERKSt6locale __gxx_personality_v0 _ZTISt9exception _ZNKSt11__use_cacheISt18__moneypunct_cacheIcLb1EEEclERKSt6locale _ZNSt16__numpunct_cacheIcEC1Em calloc _ZN5Utils4trimESs _ZNKSt10moneypunctIcLb0EE16do_thousands_sepEv _ZNKSt8numpunctIcE12do_falsenameEv _ZNKSs4rendEv _ZNSt14basic_ofstreamIcSt11char_traitsIcEE4openERKSsSt13_Ios_Openmode _ZNKSs4findERKSsm _ZTSSt15messages_bynameIcE _ZNSt8ios_base7failureD0Ev _ZNSt18__moneypunct_cacheIcLb1EED2Ev _ZNKSt11__use_cacheISt18__moneypunct_cacheIcLb0EEEclERKSt6locale malloc_usable_size __register_frame_info_bases _ZTSSt9time_base _ZNKSt11__timepunctIcE15_M_date_formatsEPPKc _ZNSt14collate_bynameIcEC1EPKcm _ZNSs6insertEmRKSs strtod _ZTISt10moneypunctIcLb1EE _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEED0Ev _ZNSdC2EPSt15basic_streambufIcSt11char_traitsIcEE _ZNSt13basic_filebufIcSt11char_traitsIcEEC2Ev _ZNSt14basic_ofstreamIcSt11char_traitsIcEED1Ev _ZNSt11regex_errorC2ENSt15regex_constants10error_typeE _ZTTSt18basic_stringstreamIcSt11char_traitsIcESaIcEE _ZNSt9type_infoD1Ev _ZN10__cxxabiv119__foreign_exceptionD1Ev _ZTSSt12domain_error write _ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEEmc _ZTISt19basic_ostringstreamIcSt11char_traitsIcESaIcEE _ZNSsC1EPKcmRKSaIcE _ZNSi10_M_extractIlEERSiRT_ _ZSt9use_facetISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZNSt8ios_base10scientificE _ZTSSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZTVSt12future_error _ZNSs4rendEv __stdio_impl_close _ZNSt9type_infoD0Ev _ZTSSt14codecvt_bynameIcc9mbstate_tE _ZNSt13runtime_errorD1Ev _ZNSt17__timepunct_cacheIcEC1Em _ZNSt13basic_filebufIcSt11char_traitsIcEE8overflowEi _ZNSt8ios_base15sync_with_stdioEb _ZNSi10_M_extractIbEERSiRT_ _ZNSi10_M_extractIfEERSiRT_ _ZNSdD2Ev fstat fprintf _ZNSs12_Alloc_hiderC2EPcRKSaIcE _ZTIN9__gnu_cxx20recursive_init_errorE _ZNSsC1ERKSsmmRKSaIcE _ZNSt12domain_errorC2ERKSs AllocMem _ZSt14__convert_to_vIeEvPKcRT_RSt12_Ios_IostateRKPi _ZNSt8ios_base11adjustfieldE _ZNSt14basic_ifstreamIcSt11char_traitsIcEED2Ev _ZNSt12domain_errorC1ERKSs _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2EiSt13_Ios_Openmodem _ZNSt12domain_errorD1Ev _ZNSsC2IPcEET_S1_RKSaIcE _ZSt9has_facetISt8numpunctIcEEbRKSt6locale _ZNSt15basic_streambufIcSt11char_traitsIcEE7pubsyncEv _ZTSSt17__timepunct_cacheIcE _ZNKSt9basic_iosIcSt11char_traitsIcEEcvPvEv _ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_ES3_RKS6_ _ZStrsIcSt11char_traitsIcESaIcEERSt13basic_istreamIT_T0_ES7_RSbIS4_S5_T1_E _ZN9__gnu_cxx15__concat_size_tEPcmm _ZTVSt16__numpunct_cacheIcE _ZNSt8ios_base4leftE _ZNSt15underflow_errorD0Ev _ZNSt14error_categoryD0Ev _ZNKSt9type_info11__do_upcastEPKN10__cxxabiv117__class_type_infoEPPv _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNSt11range_errorD2Ev _ZNSt10moneypunctIcLb1EED0Ev _ZNSolsEPFRSt8ios_baseS0_E _ZNSolsEe _ZNSs7replaceEmmPKc _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE12_M_group_intEPKcmcRSt8ios_basePcS9_Ri _ZNSaIcED1Ev _ZTVSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Em _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE24_M_extract_wday_or_monthES3_S3_RiPPKcmRSt8ios_baseRSt12_Ios_Iostate ReceiveMessageM __deregister_frame_info _ZNSo6sentryC2ERSo _ZSt13get_terminatev _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPKv _ZNSt5ctypeIcE2idE _ZTv0_n12_NSt14basic_ifstreamIcSt11char_traitsIcEED0Ev _stdout_buf _ZNSt12__basic_fileIcE8sys_openEiSt13_Ios_Openmode _ZNSt15underflow_errorC2ERKSs _ZNSs7replaceEmmRKSsmm _ZNSt15basic_streambufIcSt11char_traitsIcEE6stosscEv _ZNSt17bad_function_callD2Ev fseeko _ZNKSs2atEm _ZNSt15basic_streambufIcSt11char_traitsIcEE5sgetcEv _ZNSs6assignERKSsmm tell _ZNSt9basic_iosIcSt11char_traitsIcEE3tieEPSo _Unwind_Resume _ZNSsC1IPcEET_S1_RKSaIcE _ZNKSs7_M_iendEv _ZNSt10ctype_base5alnumE _Unwind_DeleteException _ZTCSt18basic_stringstreamIcSt11char_traitsIcESaIcEE0_Sd _ZNSt10__num_base12_S_atoms_outE fseek _ZNKSt5ctypeIcE9do_narrowEcc _ZNKSt8numpunctIcE16do_thousands_sepEv _ITM_registerTMCloneTable SendMessageM _ZNSt11__timepunctIcEC1EPiPKcm _ZNSt13basic_filebufIcSt11char_traitsIcEE16_M_destroy_pbackEv _ZNKSs5beginEv _ZNSt13basic_filebufIcSt11char_traitsIcEE7seekposESt4fposI9mbstate_tESt13_Ios_Openmode _ZTISt17moneypunct_bynameIcLb1EE _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1EP4FILESt13_Ios_Openmodem Close _ZN10__cxxabiv121__vmi_class_type_infoD2Ev _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE15_M_insert_floatIdEES3_S3_RSt8ios_baseccT_ _ZNSt8ios_base8internalE _ZTVSt15numpunct_bynameIcE _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_mc _ZNSs4_Rep20_S_empty_rep_storageE _ZNKSt10moneypunctIcLb1EE11do_groupingEv _ZNSt15basic_streambufIcSt11char_traitsIcEE5imbueERKSt6locale _ZNSo9_M_insertImEERSoT_ _ZNSi3getERSt15basic_streambufIcSt11char_traitsIcEE _ZNKSt13runtime_error4whatEv _ZNSt8ios_base3ateE _ZNKSt8messagesIcE4openERKSsRKSt6locale _ZTVSt21__ctype_abstract_baseIcE _ZTISt13runtime_error _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St13_Setprecision _ZNK10__cxxabiv117__class_type_info11__do_upcastEPKS0_PPv _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE6setbufEPcl _ZZNSt13basic_filebufIcSt11char_traitsIcEE5closeEvEN14__close_sentryD1Ev _ZNSt13basic_filebufIcSt11char_traitsIcEE6setbufEPcl _ZNSt6locale4noneE _ZNSt15basic_streambufIcSt11char_traitsIcEE9underflowEv _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intItEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ __fseeko_unlocked _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1EPKcm _ZTSSt13bad_exception _ZTSSt15numpunct_bynameIcE _ZNSt8numpunctIcE2idE _ZNKSt10moneypunctIcLb1EE16do_negative_signEv _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEED2Ev memchr _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEEC1ERKSsSt13_Ios_Openmode __fini_stdio _ZTVSt12length_error _ZNSt15basic_streambufIcSt11char_traitsIcEE12__safe_pbumpEl _ZNKSt8messagesIcE20_M_convert_from_charEPc _ZNSt10ctype_base5punctE _ZNKSt20bad_array_new_length4whatEv Exit _ZNKSt8bad_cast4whatEv _ZTISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZNSt8ios_base8showbaseE stdin _ZTISt11__timepunctIcE _ZTVSt14collate_bynameIcE _ZNKSt8messagesIcE3getEiiiRKSs _ZTISt14codecvt_bynameIcc9mbstate_tE _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecd _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_S2_S2_ _ZNKSt9basic_iosIcSt11char_traitsIcEE3tieEv _ZTISt12codecvt_base _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE4fileEv _ZNSsC1ERKSaIcE _ZNSt8ios_base7unitbufE _ZNSolsEs _ZNSt14basic_ifstreamIcSt11char_traitsIcEE5closeEv _ZN5Utils10inportByteEt _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEED2Ev _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx _ZNSs4_Rep15_M_set_sharableEv _ZTv0_n12_NSt19basic_ostringstreamIcSt11char_traitsIcESaIcEED0Ev _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basece _ZTv0_n12_NSt18basic_stringstreamIcSt11char_traitsIcESaIcEED1Ev _ZNSs4backEv _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1Ev _ZN6Logger3logEPKcPc _ZNSt8ios_base17_M_call_callbacksENS_5eventE _ZNKSt10moneypunctIcLb1EE14do_curr_symbolEv _ZNKSt5ctypeIcE2isEjc _ZNSs4_Rep11_S_max_sizeE WriteS _ZNSt16invalid_argumentD2Ev _ZNSoD0Ev _ZNSt5ctypeIcEC1EPKjbm _ZNKSt8numpunctIcE11do_truenameEv _ZNSi7getlineEPclc _ZNSt12length_errorD1Ev _ZSt9use_facetISt8messagesIcEERKT_RKSt6locale _start _ZNSt15basic_streambufIcSt11char_traitsIcEE8in_availEv _ZTISt11logic_error _ZNSt8numpunctIcED2Ev __deregister_frame_info_bases _ZNKSs4dataEv _ZNKSt7collateIcE4hashEPKcS2_ _ZNSaIwED2Ev _ZTSSt9basic_iosIcSt11char_traitsIcEE _ZNSt12__basic_fileIcE5closeEv _ZGVNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNSo5seekpESt4fposI9mbstate_tE _ZTSSt9type_info _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEEC2ERKSsSt13_Ios_Openmode _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC1EiSt13_Ios_Openmodem _ZNKSs4cendEv _ZNKSs8capacityEv _ZNSs7_M_dataEPc _ZNSt8numpunctIcED1Ev AtomicBlockDual _ZNSt15underflow_errorC1ERKSs _ZNKSt9bad_alloc4whatEv _ZNSoC1EPSt15basic_streambufIcSt11char_traitsIcEE _ZTVSt14codecvt_bynameIcc9mbstate_tE __cxa_pure_virtual _ZNSt15numpunct_bynameIcED2Ev _ZTISt16__numpunct_cacheIcE ftello _ZNKSs8_M_limitEmm __stdio_impl_fileno _ZTVSt9bad_alloc _ZNSolsEi _ZNSt7codecvtIcc9mbstate_tEC1Em _ZTVSt7collateIcE _Z13waitForBuffer11Ps2Buffer_t signal _ZNKSs7crbeginEv read _ZNSs14_M_replace_auxEmmmc _ZNSt10moneypunctIcLb0EEC1EPSt18__moneypunct_cacheIcLb0EEm _ZNSo5tellpEv _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1EPKcSt13_Ios_Openmode _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_yearES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNSsC2ERKSs _Z15handleMouseDatah _ZStorSt13_Ios_OpenmodeS_ _ZNKSs13get_allocatorEv _ZTISt10bad_typeid _ZNSt10money_base8_S_atomsE __fclose_static_unlocked _ZTVSt20bad_array_new_length _ZTSSt9bad_alloc _ZNSt13basic_fstreamIcSt11char_traitsIcEEC2ERKSsSt13_Ios_Openmode _ZNSt8ios_base9uppercaseE _ZNSt12__basic_fileIcE9showmanycEv _ZNKSt18basic_stringstreamIcSt11char_traitsIcESaIcEE5rdbufEv strcoll _ZNSt8ios_baseC2Ev isupper _ZNSt8ios_base4InitD2Ev __stdio_impl_eof _ZTISt13basic_fstreamIcSt11char_traitsIcEE _ZNSolsEx _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRd _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_a _ZNKSt10moneypunctIcLb0EE16do_negative_signEv _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEED2Ev _ZNKSi6gcountEv _ZNKSs4findEPKcmm _ZNSt15basic_streambufIcSt11char_traitsIcEE8pubimbueERKSt6locale _ZNKSt8numpunctIcE9falsenameEv _ZTCSd8_So _ZNSs5eraseEN9__gnu_cxx17__normal_iteratorIPcSsEES2_ _ZNKSt10moneypunctIcLb1EE13positive_signEv _ZN6Logger3logESsz _ZTv0_n12_NSdD1Ev _ZGVNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNSolsEj _ZTISt12system_error _ZGVNSt10moneypunctIcLb1EE2idE _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb1EEES3_S3_RSt8ios_basecRKSs _ZNSt6locale7classicEv _ZNKSt8messagesIcE18_M_convert_to_charERKSs _ZTCSt13basic_fstreamIcSt11char_traitsIcEE8_So _ZNKSt14basic_ifstreamIcSt11char_traitsIcEE5rdbufEv _ZNSt12domain_errorD2Ev strncpy _ZNKSs7compareERKSs _ZNKSt15basic_streambufIcSt11char_traitsIcEE6getlocEv _ZNKSt7codecvtIcc9mbstate_tE9do_lengthERS0_PKcS4_m _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Em __open_file_list _ZNSs7_M_leakEv __init_stdio _ZTVN10__cxxabiv119__foreign_exceptionE _ZNSt20bad_array_new_lengthD0Ev _ZNSi3getERc _ZNSt15numpunct_bynameIcED1Ev ShareMem __cxa_throw_bad_array_new_length _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC1Ev _ZNSt9type_infoD2Ev _ZNSt15basic_streambufIcSt11char_traitsIcEE10pubseekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZNKSt11__timepunctIcE6_M_putEPcmPKcPK2tm _ZN10__cxxabiv119__foreign_exceptionD0Ev _ZNSt8ios_base3decE _ZNK10__cxxabiv120__si_class_type_info11__do_upcastEPKNS_17__class_type_infoEPKvRNS1_15__upcast_resultE _ZNSt8ios_base7_M_initEv _ZNSt16invalid_argumentD1Ev _ZNKSs3endEv _ZNSoC2Ev realloc _ZTINSt6locale5facetE _ZTSN10__cxxabiv121__vmi_class_type_infoE _ZNSi4readEPcl _ZNSs9_M_assignEPcmc _ZThn8_NSt13basic_fstreamIcSt11char_traitsIcEED0Ev _ZTSSt18__moneypunct_cacheIcLb1EE _ZSt9has_facetISt5ctypeIcEEbRKSt6locale _ZGVNSt10moneypunctIcLb0EE2idE _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecb _ZNKSs5rfindEcm _ZGVNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE __cxa_atexit _ZNSaIcEC2Ev _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt5ctypeIcED1Ev _ZNSt8ios_base13_M_grow_wordsEib _ZTSSt15underflow_error _ZNSi3getERSt15basic_streambufIcSt11char_traitsIcEEc _ZTSSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE8overflowEi _ZTIN10__cxxabiv119__foreign_exceptionE _ZNKSs13find_first_ofEcm _ZNKSt11__timepunctIcE9_M_monthsEPPKc _ZNSt15messages_bynameIcED0Ev _ZNSt15underflow_errorD2Ev _ZTSSt10ctype_base _ZNSt18__moneypunct_cacheIcLb1EED1Ev _ZNSt10moneypunctIcLb1EE2idE _ZTSSd _ZNSo9_M_insertIyEERSoT_ _ZNKSt7codecvtIcc9mbstate_tE11do_encodingEv _ZTVSt8numpunctIcE _ZNKSt9basic_iosIcSt11char_traitsIcEE5widenEc _ZNSt17moneypunct_bynameIcLb0EEC2EPKcm __x86.get_pc_thunk.bx _ZNKSt8numpunctIcE11do_groupingEv _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIxEES3_S3_RSt8ios_basecT_ _ZNSt17moneypunct_bynameIcLb0EED0Ev mouseReceiverTransaction _ZNSt15basic_streambufIcSt11char_traitsIcEE7seekposESt4fposI9mbstate_tESt13_Ios_Openmode _ZNSiC1Ev memcmp _ZSt4endsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ _ZNSt10moneypunctIcLb0EE4intlE _ZNSt6localeD1Ev _ZN5Utils11outportByteEth _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St13_Setprecision _ZTVN9__gnu_cxx20recursive_init_errorE malloc_trim _ZTVSt17__timepunct_cacheIcE _ZNSt9bad_allocD0Ev fdopen _ZNKSt5ctypeIcE10do_toupperEc _ZN10__cxxabiv120__si_class_type_infoD1Ev _ZNKSt9basic_iosIcSt11char_traitsIcEE7rdstateEv _ZNSs13shrink_to_fitEv _ZNSt6locale9_S_globalE sscanf _ZNSt9basic_iosIcSt11char_traitsIcEE5rdbufEPSt15basic_streambufIcS1_E _ZNSt15basic_streambufIcSt11char_traitsIcEE4syncEv _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEEC1ESt13_Ios_Openmode _ZNSt11range_errorD1Ev _ZTSSt11range_error _Unwind_RaiseException _ZNSt7collateIcEC1Em isalpha _ZN9__gnu_cxx15__snprintf_liteEPcmPKcS0_ _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe _ZNKSt10moneypunctIcLb1EE13negative_signEv _ZTISt12domain_error _ZNKSt9type_info14__is_pointer_pEv _ZTSSt8bad_cast _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEEC1ERKSsSt13_Ios_Openmode _ZNSt10ctype_base5cntrlE _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_NS0_IPKcSsEES5_ _ZTISt8messagesIcE _ZTISt14overflow_error _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt6locale5_Impl19_M_replace_categoryEPKS0_PKPKNS_2idE _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE9_M_insertILb0EEES3_S3_RSt8ios_basecRKSs _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE17_M_stringbuf_initESt13_Ios_Openmode _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEEC1ERKSsSt13_Ios_Openmode _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St8_SetfillIS3_E _ZNSt8ios_base4InitC1Ev fread _ZTVSt9exception _ZN10__cxxabiv115__forced_unwindD0Ev _ZNSt12__basic_fileIcEC2EPi _ZNSt8ios_base9boolalphaE _ZNSt8ios_base3endE _ZTSSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_RKSs _ZNSt15basic_streambufIcSt11char_traitsIcEED2Ev _ZNSt6localeaSERKS_ CliArgsRelease _ZNK10__cxxabiv117__class_type_info20__do_find_public_srcElPKvPKS0_S2_ _ZNSs5clearEv _ITM_deregisterTMCloneTable sbrk _ZSt20__throw_domain_errorPKc _InitLibc _ZNSt6locale5ctypeE _ZSt19__throw_logic_errorPKc _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10date_orderEv _ZTVN10__cxxabiv117__class_type_infoE __cxa_throw _ZNKSs13find_first_ofEPKcmm _Unwind_SetIP _ZNKSt10moneypunctIcLb0EE13negative_signEv _ZNSt16__numpunct_cacheIcE8_M_cacheERKSt6locale _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE6xsgetnEPcl _ZNSt18basic_stringstreamIcSt11char_traitsIcESaIcEEC2ERKSsSt13_Ios_Openmode _ZNSt10moneypunctIcLb1EED1Ev _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIyEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZTISt12length_error _ZNKSs12find_last_ofEcm _ZNKSt9basic_iosIcSt11char_traitsIcEE4failEv _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St12_Setiosflags _ZNSs4_Rep13_M_set_leakedEv _ZNSt9basic_iosIcSt11char_traitsIcEE4fillEc _ZNSi10_M_extractIxEERSiRT_ _ZSt19__throw_range_errorPKc _ZNSsC2EPKcmRKSaIcE _ZNSt16invalid_argumentC1ERKSs fopen _Z21registerOperationModev __bss_start _ZNSt10moneypunctIcLb1EED2Ev _ZNKSs13find_first_ofERKSsm _ZNSt9basic_iosIcSt11char_traitsIcEEC1Ev _ZNSt8ios_base3appE AtomicBlock _ZNSt11__timepunctIcED0Ev _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEEC1ERKSsSt13_Ios_Openmode _ZTVSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZNSt6locale5facetD2Ev _ZNKSs7compareEmmRKSs memset _ZNSt15basic_streambufIcSt11char_traitsIcEE7seekoffExSt12_Ios_SeekdirSt13_Ios_Openmode _ZNSs4_Rep26_M_set_length_and_sharableEm __vfprintf_unlocked _ZNSs12_S_empty_repEv main _ZTSSt13runtime_error _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE15_M_extract_nameES3_S3_RiPPKcmRSt8ios_baseRSt12_Ios_Iostate _ZNSt7collateIcED1Ev _ZNSt13basic_fstreamIcSt11char_traitsIcEE5closeEv _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecl _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St14_Resetiosflags _ZNKSt8messagesIcE6do_getEiiiRKSs _ZNSt8messagesIcED0Ev AtomicTryLockDual _ZNSt15basic_streambufIcSt11char_traitsIcEE4setgEPcS3_S3_ _ZNSt8ios_base3hexE _ZTISt18__moneypunct_cacheIcLb0EE AtomicLock _ZTSSt15basic_streambufIcSt11char_traitsIcEE _ZTISt19basic_istringstreamIcSt11char_traitsIcESaIcEE _ZNSt15basic_streambufIcSt11char_traitsIcEEaSERKS2_ _ZTVSt10bad_typeid _ZNKSt15basic_streambufIcSt11char_traitsIcEE5epptrEv _ZNKSt10moneypunctIcLb1EE14do_frac_digitsEv _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED0Ev ftell _ZTTSd _ZNSt14basic_ofstreamIcSt11char_traitsIcEED0Ev _ZTSSt15basic_stringbufIcSt11char_traitsIcESaIcEE _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEED1Ev _ZNKSt9basic_iosIcSt11char_traitsIcEE4fillEv _ZSt21__throw_bad_exceptionv __cxa_get_globals_fast strxfrm _ZNSt6locale21_S_normalize_categoryEi parseargs _ZNSsaSEOSs _ZSt5flushIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ _ZNSt12__basic_fileIcED2Ev _stdout _ZTVSt18__moneypunct_cacheIcLb0EE GetTid _ZSt25__throw_bad_function_callv _ZN9__gnu_cxx20recursive_init_errorD0Ev _ZTSNSt8ios_base7failureE Millis _ZTVSt14error_category _ZTSSi _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEED1Ev _ZNSirsERx _ZNSt5ctypeIcED0Ev _ZTVSt8bad_cast _ZdaPv _ZNSt10moneypunctIcLb0EED1Ev mallopt _ZNKSt10bad_typeid4whatEv _ZSt13__int_to_charIcmEiPT_T0_PKS0_St13_Ios_Fmtflagsb _ZNKSt10moneypunctIcLb1EE8groupingEv _ZNSt15messages_bynameIcED1Ev fclose _ZNSt14error_categoryD1Ev _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC1ERKSsSt13_Ios_Openmode _ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Ra _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEED1Ev _ZTISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZNSt12out_of_rangeD1Ev _ZNSt8ios_base6xallocEv _ZNSt18__moneypunct_cacheIcLb0EEC2Em _ZNSt14basic_ifstreamIcSt11char_traitsIcEED1Ev _ZNSt14collate_bynameIcED2Ev _ZNKSt17bad_function_call4whatEv _ZNSsC2IPKcEET_S2_RKSaIcE _ZNSt6locale5facet15_S_get_c_localeEv time _ZNSt18__moneypunct_cacheIcLb0EED1Ev _ZNKSt8numpunctIcE16do_decimal_pointEv __stdio_impl_tell _ZNKSt13bad_exception4whatEv _ZNSspLESt16initializer_listIcE _ZNSsC2ERKSaIcE __register_frame_info_table_bases _ZSt9use_facetISt7codecvtIcc9mbstate_tEERKT_RKSt6locale _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_S1_S1_ _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE6xsputnEPKcl _ZNKSt9basic_iosIcSt11char_traitsIcEE10exceptionsEv _ZNSt14overflow_errorC2ERKSs isgraph _ZNSt11range_errorD0Ev _ZSt15future_categoryv _ZTISt17moneypunct_bynameIcLb0EE _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSt14codecvt_bynameIcc9mbstate_tEC1EPKcm _ZTSSt16bad_array_length _ZTIN10__cxxabiv117__class_type_infoE _ZNKSt14error_category23default_error_conditionEi __fflush_read_unlocked isalnum _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecy _ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE6_M_getEv _ZTCSt19basic_istringstreamIcSt11char_traitsIcESaIcEE0_Si mouseReceiverTid _ZTVSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZNSo9_M_insertIPKvEERSoT_ isprint _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSs12find_last_ofEPKcmm _ZNSt13bad_exceptionD1Ev _ZTISt20bad_array_new_length _ZNSoC1Ev _ZTVN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEE putc _ZNSt18__moneypunct_cacheIcLb0EED0Ev _ZSt9use_facetISt10moneypunctIcLb1EEERKT_RKSt6locale _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2Ev _ZNSirsERb _ZNSt13basic_fstreamIcSt11char_traitsIcEED1Ev _ZNKSt10moneypunctIcLb1EE13decimal_pointEv _ZTISt5ctypeIcE _ZNSt9basic_iosIcSt11char_traitsIcEED0Ev _ZNSoD2Ev _ZNKSt10moneypunctIcLb0EE13thousands_sepEv _ZTVSt12system_error _ZNKSt9basic_iosIcSt11char_traitsIcEE3badEv _ZNSo9_M_insertIbEERSoT_ _ZNSs6appendERKSs _ZNSs9push_backEc strcmp _ZTSSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE RegisterIrqHandler _ZNSs13_S_copy_charsEPcPKcS1_ _ZNKSt19istreambuf_iteratorIcSt11char_traitsIcEE5equalERKS2_ _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecd _ZNSt8ios_base3octE _Z15initializeMousev _ZSt4clog _ZNSt11__timepunctIcE23_M_initialize_timepunctEPi _ZNKSt7codecvtIcc9mbstate_tE13do_max_lengthEv _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC1Em _ZTVN10__cxxabiv115__forced_unwindE _ZNSi6ignoreEl _ZNSt8ios_base7failureD2Ev _ZNSt13basic_fstreamIcSt11char_traitsIcEED2Ev _ZNSt8ios_base7failureC1ERKSs _ZNSi5seekgExSt12_Ios_Seekdir _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSt11regex_errorC1ENSt15regex_constants10error_typeE _ZSt9has_facetISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZNSt10ctype_base5upperE _ZNSsC1EPKcRKSaIcE _ZNSt13basic_filebufIcSt11char_traitsIcEED1Ev _ZNSt10moneypunctIcLb0EEC1Em _ZNKSt14error_category10equivalentERKSt10error_codei _ZNSt13basic_filebufIcSt11char_traitsIcEE7_M_seekExSt12_Ios_Seekdir9mbstate_t _ZNSt8bad_castD2Ev __deregister_frame _ZNSt12out_of_rangeC1ERKSs _ZNSt11__timepunctIcE2idE malloc_footprint _fini _ZTISt18basic_stringstreamIcSt11char_traitsIcESaIcEE _ZNSt8ios_baseD0Ev _ZNSt15numpunct_bynameIcEC1EPKcm _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE8_M_pbumpEPcS4_x _ZNSs12_S_constructIPcEES0_T_S1_RKSaIcESt20forward_iterator_tag _ZTv0_n12_NSt18basic_stringstreamIcSt11char_traitsIcESaIcEED0Ev _ZN10__cxxabiv120__si_class_type_infoD0Ev _ZNSs6insertEmPKc _ZNKSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_bRSt8ios_basecRKSs _ZNSs8pop_backEv _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb0EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs _ZStrsIcSt11char_traitsIcEERSt13basic_istreamIT_T0_ES6_St5_Setw _ZTIN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE AtomicLockDual malloc_set_footprint_limit _ZNSt15basic_streambufIcSt11char_traitsIcEE5sputcEc memalign _ZTISt13basic_filebufIcSt11char_traitsIcEE sprintf _ZNSt11__timepunctIcEC1EPSt17__timepunct_cacheIcEm _ZNSt11logic_errorD2Ev _ZNSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSi5tellgEv _ZNSt16__numpunct_cacheIcEC2Em _ZNSs12_M_leak_hardEv _ZN9__gnu_cxx4ropeIcSaIcEE8_S_fetchEPNS_13_Rope_RopeRepIcS1_EEm _ZNSt10moneypunctIcLb1EEC1Em _ZTVSt17moneypunct_bynameIcLb1EE _ZTVSt10moneypunctIcLb0EE _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE15_M_insert_floatIeEES3_S3_RSt8ios_baseccT_ _ZTSSt11logic_error _ZTv0_n12_NSt19basic_ostringstreamIcSt11char_traitsIcESaIcEED1Ev _ZNSt11logic_errorD1Ev strtof _ZNSt16bad_array_lengthD0Ev _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRt _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Em _ZNSt6localeD2Ev _ZTISt11range_error _ZNSolsEPFRSt9basic_iosIcSt11char_traitsIcEES3_E __cxa_guard_release _ZNKSt8numpunctIcE13decimal_pointEv _ZNSt11range_errorC1ERKSs _ZTISt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_numES3_S3_RiiimRSt8ios_baseRSt12_Ios_Iostate _ZNKSt14error_category10equivalentEiRKSt15error_condition _ZTv0_n12_NSt19basic_istringstreamIcSt11char_traitsIcESaIcEED1Ev _Z18handleKeyboardDatah _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm __cxa_bad_cast _ZTv0_n12_NSdD0Ev _ZNSt12out_of_rangeD0Ev setlocale _ZSt3cin _ZTSSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZNSiC2Ev _ZNSiD1Ev _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE9underflowEv _Unwind_GetTextRelBase _ZTSN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEE _ZTVN10__cxxabiv121__vmi_class_type_infoE _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe __cxa_call_terminate _ZNSt6locale7numericE stderr _ZNSt8ios_base9basefieldE _ZNSt10moneypunctIcLb0EEC2EPiPKcm _ZSt9use_facetISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale __setdefbuf_unlocked _ZTIN10__cxxabiv115__forced_unwindE _ZNSo8_M_writeEPKcl __open_file_list_add _ZNKSt19basic_istringstreamIcSt11char_traitsIcESaIcEE5rdbufEv _ZNSt6locale8messagesE _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEED2Ev _ZTSSt13messages_base _ZTTSi _ZNSt15basic_streambufIcSt11char_traitsIcEEC2ERKS2_ _ZNSt5ctypeIcED2Ev _ZSt9use_facetISt7collateIcEERKT_RKSt6locale _ZNSt11regex_errorD2Ev _ZTISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZTISt17__timepunct_cacheIcE _ZTISt12future_error _ZNSi10_M_extractIyEERSiRT_ _ZSt9has_facetISt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZNSt14collate_bynameIcED0Ev _ZStplIcSt11char_traitsIcESaIcEESbIT_T0_T1_ERKS6_S8_ _ZNSt8ios_base7goodbitE _ZNSt10moneypunctIcLb1EE24_M_initialize_moneypunctEPiPKc _ZSt9has_facetISt7collateIcEEbRKSt6locale _ZNSt14codecvt_bynameIcc9mbstate_tED0Ev _ZSt14get_unexpectedv _ZNSt8ios_base4InitD1Ev _ZNKSs8_M_checkEmPKc _ZNKSs17find_first_not_ofEPKcm _ZNSt6locale5_Impl10_S_id_timeE _ZNSt10moneypunctIcLb1EEC2EPiPKcm _ZNSt8ios_base2inE _ZNKSs5emptyEv _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecx _Unwind_FindEnclosingFunction _ZN9__gnu_cxxeqIPcSsEEbRKNS_17__normal_iteratorIT_T0_EES7_ valloc _ZNSaIwEC1ERKS_ ReceiveMessageT _ZTVSt15basic_stringbufIcSt11char_traitsIcESaIcEE RegisterSignalHandler _ZTv0_n12_NSiD1Ev _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEED0Ev fputc _ZTISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE _ZTVSt5ctypeIcE _ZNSt12__basic_fileIcE8sys_openEP4FILESt13_Ios_Openmode _Znam __stdio_impl_seek __parse_mode_flags _ZNSs5eraseEmm _ZNKSt11__timepunctIcE15_M_am_pm_formatEPKc _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRl _ZTSN10__cxxabiv119__foreign_exceptionE _ZNKSs5rfindERKSsm _ZNSdC2Ev _ZNSi6sentryC1ERSib _ZNSsC2ERKSsmm mallinfo _ZNKSs16find_last_not_ofERKSsm _ZSt9has_facetISt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEEbRKSt6locale _ZNKSt7collateIcE7do_hashEPKcS2_ _ZNSt6locale5_ImplC1ERKS0_m _ZTVSt15basic_streambufIcSt11char_traitsIcEE _ZNKSt10moneypunctIcLb1EE16do_decimal_pointEv _ZNKSt5ctypeIcE9do_narrowEPKcS2_cPc _ZNSt12system_errorD0Ev __fclose_static _ZNSt12future_errorD2Ev _ZNSt16bad_array_lengthD1Ev _Unwind_GetLanguageSpecificData _ZTISt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE __cxa_guard_abort ReceiveMessageTM _ZNSt10moneypunctIcLb1EEC1EPSt18__moneypunct_cacheIcLb1EEm _ZNSt16invalid_argumentD0Ev _ZNSt13basic_fstreamIcSt11char_traitsIcEEC1ERKSsSt13_Ios_Openmode _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEEC2ERKSsSt13_Ios_Openmode _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE9pbackfailEi _ZTCSt18basic_stringstreamIcSt11char_traitsIcESaIcEE0_Si _ZNSt15basic_streambufIcSt11char_traitsIcEE9sputbackcEc sharedArea _ZNSt8ios_baseD2Ev __cxa_begin_catch _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED1Ev _ZNSs6assignESt16initializer_listIcE _ZNSt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZN10__cxxabiv117__class_type_infoD2Ev _ZNSt6locale5facet9_S_c_nameE _ZN10__cxxabiv112__unexpectedEPFvvE _ZNSsC2EOSs _ZNSt9basic_iosIcSt11char_traitsIcEE10exceptionsESt12_Ios_Iostate _ZNKSt10moneypunctIcLb0EE11curr_symbolEv _ZNSt17bad_function_callD0Ev _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode _ZThn8_NSt18basic_stringstreamIcSt11char_traitsIcESaIcEED0Ev _ZTSSt12length_error _ZNKSt11__timepunctIcE20_M_date_time_formatsEPPKc OpenFS _ZNSt13basic_fstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode strftime _ZTSSt17bad_function_call _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14do_get_weekdayES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNSi10_M_extractIjEERSiRT_ _ZNSt17bad_function_callD1Ev kvlog _ZStlsISt11char_traitsIcEERSt13basic_ostreamIcT_ES5_PKa _ZNSt14basic_ofstreamIcSt11char_traitsIcEEC2ERKSsSt13_Ios_Openmode _ZSt16__throw_bad_castv _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIjEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZNKSt8numpunctIcE8truenameEv __fdopen_static __ftello_unlocked _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2EP4FILESt13_Ios_Openmodem _ZNSt13bad_exceptionD0Ev _ZTSSt14basic_ofstreamIcSt11char_traitsIcEE _ZNSt14basic_ofstreamIcSt11char_traitsIcEE5closeEv _ZN10__cxxabiv119__terminate_handlerE __gcclibcxx_demangle_callback _ZNSt11__timepunctIcED1Ev _ZNSo5seekpExSt12_Ios_Seekdir _ZTVSt15underflow_error _ZNKSt18basic_stringstreamIcSt11char_traitsIcESaIcEE3strEv _ZNSt13basic_filebufIcSt11char_traitsIcEE22_M_convert_to_externalEPcl _ZNSt6locale8monetaryE _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2ERKSsSt13_Ios_Openmode _ZNK10__cxxabiv121__vmi_class_type_info12__do_dyncastElNS_17__class_type_info10__sub_kindEPKS1_PKvS4_S6_RNS1_16__dyncast_resultE _ZNKSt8numpunctIcE13thousands_sepEv _ZSt9use_facetISt5ctypeIcEERKT_RKSt6locale _ZNSs10_S_compareEmm _ZNSt8ios_base4Init11_S_refcountE _ZNKSo6sentrycvbEv _ZNSt6locale5_Impl13_S_id_collateE __cxa_allocate_exception _ZNKSt11__timepunctIcE21_M_months_abbreviatedEPPKc _ZNKSt19basic_istringstreamIcSt11char_traitsIcESaIcEE3strEv fwrite _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRe _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecl _ZNSt11regex_errorD0Ev _ZNKSt14basic_ofstreamIcSt11char_traitsIcEE5rdbufEv _ZN14__gnu_internal8buf_coutE _ZNSt13basic_filebufIcSt11char_traitsIcEE13_M_set_bufferEl _ZNSt18__moneypunct_cacheIcLb0EED2Ev _ZTIN10__cxxabiv120__si_class_type_infoE _ZNKSt7codecvtIcc9mbstate_tE5do_inERS0_PKcS4_RS4_PcS6_RS6_ _ZNSo6sentryC1ERSo _ZNKSt12__basic_fileIcE7is_openEv _ZNSt17__timepunct_cacheIcED2Ev _ZSt15set_new_handlerPFvvE _ZNSirsERl _ZNSsaSEc _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEC1Em SetWorkingDirectoryP _Unwind_ForcedUnwind _ZNSt13basic_filebufIcSt11char_traitsIcEED2Ev _edata _ZNKSi6sentrycvbEv packetsCount _ZNSt5ctypeIcE13classic_tableEv _ZNKSt10moneypunctIcLb0EE13do_pos_formatEv _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRy _ZNSt15basic_streambufIcSt11char_traitsIcEE6snextcEv _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE7seekposESt4fposI9mbstate_tESt13_Ios_Openmode _ZTVSt9basic_iosIcSt11char_traitsIcEE _ZNSi10_M_extractIPvEERSiRT_ _ZNSt6locale5facet18_S_create_c_localeERPiPKcS1_ _end _ZSt7nothrow _ZNSiD2Ev _ZNSt8ios_base3curE _ZNSt13runtime_errorD0Ev _ZNSirsEPFRSt8ios_baseS0_E mousePacketBuffer _ZNSt13basic_filebufIcSt11char_traitsIcEE26_M_destroy_internal_bufferEv _ZNSs4_Rep8_M_cloneERKSaIcEm _ZTVSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE6do_putES3_RSt8ios_basecPK2tmcc _ZNSt15basic_streambufIcSt11char_traitsIcEE10pubseekposESt4fposI9mbstate_tESt13_Ios_Openmode _ZNSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED0Ev _ZNSsC1EOSs __RestoreInterruptedStateCallback _ZSt9has_facetISt11__timepunctIcEEbRKSt6locale _ZTSSt11__timepunctIcE _ZSt4endlIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_ _ZNSirsERe _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEED0Ev _ZNKSs6cbeginEv _ZThn8_NSt13basic_fstreamIcSt11char_traitsIcEED1Ev _ZNKSt5ctypeIcE8do_widenEc _ZNSaIcEC1ERKS_ _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16_M_extract_floatES3_S3_RSt8ios_baseRSt12_Ios_IostateRSs _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEED1Ev __ExitThread _ZNSt15basic_streambufIcSt11char_traitsIcEE7sungetcEv _ZNSi8readsomeEPcl _ZTv0_n12_NSoD1Ev _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEE3strERKSs _ZNK10__cxxabiv117__class_type_info12__do_dyncastElNS0_10__sub_kindEPKS0_PKvS3_S5_RNS0_16__dyncast_resultE _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_bRSt8ios_baseRSt12_Ios_IostateRe _ZSt21__copy_streambufs_eofIcSt11char_traitsIcEElPSt15basic_streambufIT_T0_ES6_Rb _ZNSt9exceptionD1Ev _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEEC1EP4FILE _ZNSt9basic_iosIcSt11char_traitsIcEEC2EPSt15basic_streambufIcS1_E _ZNSt10moneypunctIcLb1EEC2EPSt18__moneypunct_cacheIcLb1EEm _ZTINSt8ios_base7failureE _ZSt4cout _ZNKSt10moneypunctIcLb0EE8groupingEv _ZNSt9basic_iosIcSt11char_traitsIcEE8setstateESt12_Ios_Iostate _ZNSt13basic_filebufIcSt11char_traitsIcEE6xsgetnEPcl _ZNSsaSESt16initializer_listIcE _ZNKSt10moneypunctIcLb1EE10neg_formatEv _ZNSt6locale7collateE _ZNKSt8time_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecPK2tmcc _ZNSi4syncEv _ZNSt6locale2id11_S_refcountE _ZTISt14basic_ifstreamIcSt11char_traitsIcEE _ZNSt11__timepunctIcEC2EPiPKcm _ZNSs4_Rep9_S_createEmmRKSaIcE _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St8_SetfillIS3_E GetExecutablePath exit _Unwind_SetGR _ZNSt8ios_base5fixedE _ZNSspLERKSs _ZTSN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEE _ZGVNSt8numpunctIcE2idE _ZNKSt12future_error4whatEv _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE6do_getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIyEES3_S3_RSt8ios_basecT_ _ZTVSt12domain_error keyboardReceiverTransaction _ZNSt14error_categoryD2Ev _ZSt9has_facetISt8messagesIcEEbRKSt6locale _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE8get_dateES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNSt15basic_streambufIcSt11char_traitsIcEE4setpEPcS3_ _ZNSt8messagesIcEC1EPiPKcm _ZNSt12__basic_fileIcE4syncEv _ZN10__cxxabiv111__terminateEPFvvE _ZNSs7replaceEmmmc _ZNSs5frontEv _ZNSt8numpunctIcEC1EPSt16__numpunct_cacheIcEm Seek _ZTVSt19basic_istringstreamIcSt11char_traitsIcESaIcEE _ZNSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEED2Ev _ZNSt12__basic_fileIcE6xsputnEPKcl _ZTISt14basic_ofstreamIcSt11char_traitsIcEE _ZNSt9bad_allocD1Ev _ZTv0_n12_NSt14basic_ifstreamIcSt11char_traitsIcEED1Ev _ZN9__gnu_cxx26__throw_insufficient_spaceEPKcS1_ _ZNK10__cxxabiv120__si_class_type_info12__do_dyncastElNS_17__class_type_info10__sub_kindEPKS1_PKvS4_S6_RNS1_16__dyncast_resultE _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE13do_date_orderEv _ZNSt5__padIcSt11char_traitsIcEE6_S_padERSt8ios_basecPcPKcll _ZTISt7collateIcE _ZNSt6locale5_Impl14_S_id_messagesE _ZTISt13bad_exception _ZTv0_n12_NSt19basic_istringstreamIcSt11char_traitsIcESaIcEED0Ev _ZTSSt21__ctype_abstract_baseIcE __open_file_list_unlock _ZNKSt9basic_iosIcSt11char_traitsIcEE4goodEv _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE9showmanycEv _ZNKSt15basic_streambufIcSt11char_traitsIcEE4pptrEv _ZNSt17moneypunct_bynameIcLb0EED1Ev _ZTISt16bad_array_length _ZNSt15time_put_bynameIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEC2EPKcm _ZTISt14collate_bynameIcE _ZNSt7codecvtIcc9mbstate_tEC2Em _ZNSt11__timepunctIcEC2EPSt17__timepunct_cacheIcEm _ZNKSt6locale2id5_M_idEv iscntrl _ZSt7setfillIcESt8_SetfillIT_ES1_ _ZNKSt5ctypeIcE14_M_narrow_initEv _ZNKSt10moneypunctIcLb0EE11frac_digitsEv _ZNSo9_M_insertIlEERSoT_ _ZNSt8ios_base5truncE _ZNSt13basic_filebufIcSt11char_traitsIcEE9underflowEv _ZNSt8messagesIcEC2EPiPKcm _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEEC2Ev _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRj _ZTVSt14basic_ofstreamIcSt11char_traitsIcEE __fflush_write_unlocked _ZNSt12domain_errorD0Ev _ZNKSt8messagesIcE7do_openERKSsRKSt6locale _ZNSt9basic_iosIcSt11char_traitsIcEED1Ev _ZNSdC1EPSt15basic_streambufIcSt11char_traitsIcEE fileno _ZNSirsERPv _ZNKSs5c_strEv _ZNSt7codecvtIcc9mbstate_tED1Ev _ZNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNSt7collateIcE2idE _ZNSt10moneypunctIcLb0EEC2EPSt18__moneypunct_cacheIcLb0EEm _ZN9__gnu_cxx18stdio_sync_filebufIcSt11char_traitsIcEE5uflowEv _ZNK10__cxxabiv121__vmi_class_type_info20__do_find_public_srcElPKvPKNS_17__class_type_infoES2_ _ZNSt14basic_ifstreamIcSt11char_traitsIcEED0Ev _ZNSt6locale13_S_categoriesE _ZNSt8ios_base7failureC2ERKSs _ZTISt10moneypunctIcLb0EE _ZNSt9basic_iosIcSt11char_traitsIcEE5clearESt12_Ios_Iostate _stderr_buf _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEEC2ESt13_Ios_Openmode _ZNSolsEd _ZSt20__throw_out_of_rangePKc _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEE2fdEv _ZNSt7codecvtIcc9mbstate_tE2idE _ZNKSs7compareEmmPKcm _ZNSs6insertEN9__gnu_cxx17__normal_iteratorIPcSsEEc _ZTVSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZNSt10moneypunctIcLb0EED0Ev _ZNSt11__timepunctIcEC1Em _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEE3strERKSs _ZNSt8ios_base4Init20_S_synced_with_stdioE _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE13_M_insert_intIlEES3_S3_RSt8ios_basecT_ _ZNSo9_M_insertIdEERSoT_ _Unwind_GetGR __cxa_get_globals _ZNSt13basic_fstreamIcSt11char_traitsIcEE4openERKSsSt13_Ios_Openmode TellS _ZNKSt15basic_streambufIcSt11char_traitsIcEE4gptrEv _ZN10__cxxabiv120__unexpected_handlerE _ZNSt8numpunctIcEC2EPim _ZNSt19basic_istringstreamIcSt11char_traitsIcESaIcEEC1ESt13_Ios_Openmode _ZNSspLEPKc _ZNSs6appendESt16initializer_listIcE _ZNKSt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE10_M_extractILb1EEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRSs _ZTISt7codecvtIcc9mbstate_tE strlen _ZNSt19basic_ostringstreamIcSt11char_traitsIcESaIcEEC1ESt13_Ios_Openmode _ZSt23__throw_underflow_errorPKc _ZTISt9type_info open _ZNSs4_Rep12_S_empty_repEv _ZNSs12_Alloc_hiderC1EPcRKSaIcE SendMessageTM toupper _ZNSt14basic_ofstreamIcSt11char_traitsIcEED2Ev _ZNSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE11do_get_timeES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZNKSt10moneypunctIcLb1EE13do_neg_formatEv _ZTSSt9exception _ZTVSt13runtime_error _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIxEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZTCSt14basic_ifstreamIcSt11char_traitsIcEE0_Si _ZN14__gnu_internal13buf_cout_syncE _ZTSSt10bad_typeid _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRPv _ZNKSs6lengthEv _ZNSt15time_get_bynameIcSt19istreambuf_iteratorIcSt11char_traitsIcEEED2Ev sig_handler_SIG_INT _ZNSs13_S_copy_charsEPcS_S_ __open_file_list_lock _ZNKSt11logic_error4whatEv _ZN5Utils10outportIntEtj _ZTSSt13basic_fstreamIcSt11char_traitsIcEE _ZNSdD0Ev __cxa_current_exception_type __fflush_unlocked _ZNSs12_S_constructIPKcEEPcT_S3_RKSaIcESt20forward_iterator_tag __cxa_bad_typeid _ZNSt9exceptionD0Ev _ZNKSt10moneypunctIcLb0EE11do_groupingEv _ZTTSt13basic_fstreamIcSt11char_traitsIcEE _ZTSSt11regex_error _ZStrsISt11char_traitsIcEERSt13basic_istreamIcT_ES5_Ph _ZTSSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE _ZNSs6resizeEmc _ZNSt15numpunct_bynameIcEC2EPKcm _ZNSt6localeC2Ev _ZNSt8numpunctIcEC1EPim _ZSt16__ostream_insertIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_PKS3_l _ZTVNSt8ios_base7failureE _ZTSSt5ctypeIcE _ZNKSt16bad_array_length4whatEv _ZN9__gnu_cxx13stdio_filebufIcSt11char_traitsIcEED1Ev _ZNSt10bad_typeidD1Ev _ZTSN9__gnu_cxx20recursive_init_errorE _ZNSt5ctypeIcE10table_sizeE _ZNSt16bad_array_lengthD2Ev fputs _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE15_M_update_egptrEv _Unwind_GetDataRelBase _ZNKSt13basic_fstreamIcSt11char_traitsIcEE5rdbufEv _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_PKcS4_ independent_comalloc _ZNSt6locale5facet11_S_c_localeE _ZNSt6locale6globalERKS_ _ZNSs6insertEmPKcm _ZNKSt14basic_ifstreamIcSt11char_traitsIcEE7is_openEv _ZNKSt9basic_iosIcSt11char_traitsIcEEntEv _ZGVNSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE2idE Log _ZNSoC2EPSt15basic_streambufIcSt11char_traitsIcEE _ZNKSt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE16do_get_monthnameES3_S3_RSt8ios_baseRSt12_Ios_IostateP2tm _ZTv0_n12_NSt13basic_fstreamIcSt11char_traitsIcEED0Ev _ZNSaIwEC2ERKS_ _ZNKSs8max_sizeEv ReadS _ZNSt6localeC1EPNS_5_ImplE _Jv_RegisterClasses _ZNSt8ios_base7failureD1Ev _ZSt9use_facetISt9money_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZTSSt17moneypunct_bynameIcLb1EE _ZNSt15basic_stringbufIcSt11char_traitsIcESaIcEE7_M_syncEPcmm _ZNSt10bad_typeidD2Ev __fwrite_unlocked _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRm _ZStlsIcSt11char_traitsIcEERSt13basic_ostreamIT_T0_ES6_St12_Setiosflags _ZNSt9basic_iosIcSt11char_traitsIcEE15_M_cache_localeERKSt6locale _ZNSt6localeC2ERKS_ _ZNSt5ctypeIcEC2EPiPKjbm _ZStlsIcSt11char_traitsIcESaIcEERSt13basic_ostreamIT_T0_ES7_RKSbIS4_S5_T1_E _ZNSs4_Rep10_M_destroyERKSaIcE _ZNKSs7compareEmmRKSsmm _ZThn8_NSdD1Ev _ZNKSs12find_last_ofERKSsm _ZNKSt10moneypunctIcLb0EE14do_frac_digitsEv _ZNSsC2EPKcRKSaIcE _ZSt7getlineIcSt11char_traitsIcESaIcEERSt13basic_istreamIT_T0_ES7_RSbIS4_S5_T1_E _ZNSt14basic_ifstreamIcSt11char_traitsIcEEC2EPKcSt13_Ios_Openmode _ZNSt8numpunctIcE22_M_initialize_numpunctEPi _ZNSs4_Rep10_M_refdataEv sched_yield _ZNSirsERs _ZTv0_n12_NSiD0Ev _ZNSs6insertEmmc _ZNSs6rbeginEv _ZN14__gnu_internal12buf_cin_syncE _ZNSiC1EPSt15basic_streambufIcSt11char_traitsIcEE _ZNKSt8messagesIcE5closeEi _ZNSt8ios_baseC1Ev __register_frame_info_table _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecy _ZNSt7codecvtIcc9mbstate_tED2Ev _Z19get_executable_namev _ZTISt13messages_base _ZTv0_n12_NSoD0Ev _ZNKSt7num_putIcSt19ostreambuf_iteratorIcSt11char_traitsIcEEE3putES3_RSt8ios_basecm _ZNSt8ios_base5rightE _ZNSt7collateIcEC2Em _ZTISt16invalid_argument _ZNKSt7collateIcE12_M_transformEPcPKcm __cxa_guard_acquire posix_memalign __register_frame_info _ZNSt17__timepunct_cacheIcED0Ev _ZNSsC2IN9__gnu_cxx17__normal_iteratorIPcSsEEEET_S4_RKSaIcE _ZNSt8numpunctIcEC2Em __stdio_impl_write _ZNSt17__timepunct_cacheIcED1Ev _ZNKSs11_M_disjunctEPKc klog _ZNSt13basic_filebufIcSt11char_traitsIcEE9pbackfailEi _ZTSSt10moneypunctIcLb0EE close _ZNSs4swapERSs _ZNSt8messagesIcED2Ev _ZNSt17moneypunct_bynameIcLb1EEC1EPKcm _ZNSt18__moneypunct_cacheIcLb1EEC1Em _ZNSt7collateIcEC2EPim _ZNSsC1EmcRKSaIcE _ZTISt14error_category _ZNSt18__moneypunct_cacheIcLb1EE8_M_cacheERKSt6locale _ZNSt13basic_filebufIcSt11char_traitsIcEED0Ev _ZNKSt10moneypunctIcLb0EE16do_positive_signEv _ZTISt8numpunctIcE _ZNSs7replaceEN9__gnu_cxx17__normal_iteratorIPcSsEES2_St16initializer_listIcE _ZTISt9money_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE __dynamic_cast _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE14_M_extract_intIlEES3_S3_S3_RSt8ios_baseRSt12_Ios_IostateRT_ _ZTSN10__cxxabiv115__forced_unwindE _ZNSt11logic_errorC1ERKSs _ZSt9use_facetISt8time_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEEERKT_RKSt6locale _ZSt20__throw_system_errori _ZNSirsERy _ZNSsC1Ev vfprintf _ZNKSt9type_info10__do_catchEPKS_PPvj _ZTSSt7codecvtIcc9mbstate_tE _ZSt14__convert_to_vIdEvPKcRT_RSt12_Ios_IostateRKPi _ZN9__gnu_cxx20recursive_init_errorD2Ev _ZNKSt9basic_iosIcSt11char_traitsIcEE5rdbufEv _ZNSt15basic_streambufIcSt11char_traitsIcEEC2Ev _ZTISi _ZNSt16invalid_argumentC2ERKSs free _ZNSt15basic_streambufIcSt11char_traitsIcEE5uflowEv _ZN9__gnu_cxx27__verbose_terminate_handlerEv _ZNKSt7num_getIcSt19istreambuf_iteratorIcSt11char_traitsIcEEE3getES3_S3_RSt8ios_baseRSt12_Ios_IostateRx _ZNSt12length_errorC2ERKSs _ZN10__cxxabiv117__class_type_infoD0Ev _ZThn8_NSt18basic_stringstreamIcSt11char_traitsIcESaIcEED1Ev __fputc_unlocked malloc_max_footprint _ZNSi3getEv _ZNSs6appendEPKcm _ZNSt13runtime_errorC1ERKSs _ZNSt14basic_ifstreamIcSt11char_traitsIcEE4openERKSsSt13_Ios_Openmode _ZNSsC1ERKSsmm 